//: version "2.1"
//: property encoding = "utf-8"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "PANIC.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"
//: require "coke"
//: require "74xxGateLevel"
//: require "tty"
//: require "m68xx"
//: require "timer"
//: require "74xx"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
supply0 w59;    //: /sn:0 {0}(211,25)(211,-12)(164,-12)(164,-1){1}
reg [7:0] w62;    //: /sn:0 {0}(#:891,749)(891,760)(701,760)(701,765){1}
reg w0;    //: /sn:0 {0}(656,208)(589,208)(589,201)(581,201){1}
//: {2}(579,199)(579,55)(390,55){3}
//: {4}(388,53)(388,-7){5}
//: {6}(388,-11)(388,-64)(378,-64){7}
//: {8}(386,-9)(338,-9)(338,-52)(-102,-52)(-102,294)(201,294){9}
//: {10}(388,57)(388,80)(389,80)(389,105){11}
//: {12}(579,203)(579,215){13}
//: {14}(581,217)(610,217)(610,1099)(547,1099){15}
//: {16}(579,219)(579,290){17}
reg w54;    //: /sn:0 {0}(234,232)(244,232)(244,217)(190,217)(190,194){1}
//: {2}(192,192)(211,192)(211,184)(635,184)(635,163)(656,163){3}
//: {4}(190,190)(190,142)(212,142){5}
//: {6}(188,192)(181,192)(181,193)(120,193){7}
reg [7:0] w8;    //: /sn:0 {0}(#:678,861)(647,861)(647,869){1}
reg [15:0] w52;    //: /sn:0 {0}(#:1187,320)(1187,469)(#:1270,469){1}
reg [15:0] w11;    //: /sn:0 {0}(#:328,1285)(328,1295)(262,1295)(262,1258)(229,1258)(#:229,1273){1}
wire [1:0] w13;    //: /sn:0 {0}(#:417,741)(417,751)(525,751){1}
//: {2}(527,749)(527,736)(428,736)(#:428,696){3}
//: {4}(527,753)(527,794){5}
wire w16;    //: /sn:0 {0}(162,1129)(167,1129)(167,1128)(191,1128){1}
//: {2}(195,1128)(218,1128)(218,1121){3}
//: {4}(220,1119)(254,1119){5}
//: {6}(218,1117)(218,1046)(771,1046)(771,988)(761,988){7}
//: {8}(193,1126)(193,1100){9}
wire [15:0] w6;    //: /sn:0 {0}(#:419,429)(419,454)(407,454)(407,477){1}
//: {2}(409,479)(564,479)(564,446){3}
//: {4}(405,479)(197,479)(197,551)(#:208,551){5}
wire w58;    //: /sn:0 {0}(673,672)(701,672)(701,718)(73,718)(73,341){1}
//: {2}(75,339)(84,339)(84,190)(99,190){3}
//: {4}(71,339)(42,339)(42,314){5}
wire w7;    //: /sn:0 {0}(458,423)(536,423)(536,422)(636,422){1}
//: {2}(640,422)(687,422)(687,406){3}
//: {4}(689,404)(702,404)(702,257){5}
//: {6}(687,402)(687,377){7}
//: {8}(638,424)(638,454)(-218,454)(-218,1187)(14,1187)(14,1174)(28,1174){9}
wire [15:0] w34;    //: /sn:0 {0}(#:473,1331)(473,1325)(472,1325)(472,1307){1}
//: {2}(#:474,1305)(686,1305)(686,1292){3}
//: {4}(472,1303)(472,1257)(505,1257)(#:505,1236){5}
wire w50;    //: /sn:0 {0}(65,934)(65,945)(35,945){1}
//: {2}(33,943)(33,868){3}
//: {4}(33,947)(33,1133)(23,1133){5}
//: {6}(19,1133)(-11,1133)(-11,1294){7}
//: {8}(-9,1296)(34,1296)(34,1287){9}
//: {10}(-11,1298)(-11,1369)(348,1369){11}
//: {12}(21,1135)(21,1169)(28,1169){13}
wire w39;    //: /sn:0 {0}(488,1400)(488,1396)(464,1396)(464,1386){1}
wire [15:0] w25;    //: /sn:0 {0}(#:404,1049)(404,1043)(412,1043)(412,1035){1}
//: {2}(412,1031)(412,988)(638,988)(638,1056)(#:646,1056){3}
//: {4}(#:410,1033)(352,1033)(352,998){5}
wire [7:0] w4;    //: /sn:0 {0}(#:391,272)(391,265){1}
//: {2}(#:393,263)(432,263)(432,248){3}
//: {4}(391,261)(391,220)(392,220)(#:392,181){5}
wire w56;    //: /sn:0 {0}(149,1152)(149,1162)(156,1162)(156,1006)(-11,1006){1}
//: {2}(-13,1004)(-13,958)(742,958)(742,744){3}
//: {4}(-13,1008)(-13,1106)(59,1106){5}
//: {6}(61,1104)(61,1065)(81,1065)(81,1096){7}
//: {8}(61,1108)(61,1119)(133,1119){9}
wire [15:0] w36;    //: /sn:0 {0}(#:383,1457)(383,1441){1}
//: {2}(383,1437)(383,1417)(384,1417)(#:384,1386){3}
//: {4}(#:381,1439)(224,1439)(224,1406){5}
wire [15:0] w22;    //: /sn:0 {0}(#:391,330)(391,336)(407,336)(407,379){1}
//: {2}(#:409,381)(532,381)(532,354){3}
//: {4}(407,383)(407,396)(419,396)(#:419,408){5}
wire w20;    //: /sn:0 {0}(673,626)(863,626)(863,654)(1053,654){1}
//: {2}(1057,654)(1059,654)(1059,597)(1088,597)(1088,578){3}
//: {4}(1055,652)(1055,433)(-254,433)(-254,679)(-321,679)(-321,724){5}
wire w60;    //: /sn:0 {0}(162,23)(181,23)(181,41)(198,41){1}
wire w29;    //: /sn:0 {0}(673,544)(734,544)(734,540)(740,540){1}
//: {2}(742,538)(742,525){3}
//: {4}(742,542)(742,723){5}
wire w30;    //: /sn:0 {0}(72,862)(377,862)(377,837){1}
//: {2}(379,835)(572,835){3}
//: {4}(576,835)(754,835){5}
//: {6}(756,833)(756,759){7}
//: {8}(758,757)(788,757)(788,747){9}
//: {10}(790,745)(800,745)(800,553)(981,553)(981,538)(971,538){11}
//: {12}(788,743)(788,738)(781,738){13}
//: {14}(756,755)(756,515){15}
//: {16}(758,513)(779,513)(779,446)(1708,446)(1708,632)(1876,632)(1876,646)(1905,646)(1905,672)(1869,672){17}
//: {18}(756,511)(756,407){19}
//: {20}(758,405)(776,405)(776,378){21}
//: {22}(754,405)(744,405){23}
//: {24}(742,403)(742,272)(752,272)(752,257){25}
//: {26}(742,407)(742,499)(125,499)(125,613){27}
//: {28}(127,615)(151,615)(151,598){29}
//: {30}(125,617)(125,652)(208,652){31}
//: {32}(756,837)(756,926)(690,926){33}
//: {34}(574,833)(574,809)(566,809){35}
//: {36}(377,833)(377,810)(369,810){37}
//: {38}(375,835)(146,835)(146,776)(150,776){39}
//: {40}(154,776)(177,776)(177,761)(165,761){41}
//: {42}(152,774)(152,769)(-47,769)(-47,739)(-282,739){43}
wire [15:0] w42;    //: /sn:0 {0}(#:770,959)(770,1001){1}
//: {2}(772,1003)(1961,1003)(1961,63){3}
//: {4}(1961,62)(1961,36){5}
//: {6}(770,1005)(770,1006)(691,1006){7}
//: {8}(687,1006)(677,1006)(677,994)(651,994)(#:651,932){9}
//: {10}(689,1008)(689,1046)(#:675,1046){11}
wire [1:0] w37;    //: /sn:0 {0}(#:50:238,696)(238,740)(152,740)(152,708)(142,708){1}
//: {2}(140,706)(#:140,681){3}
//: {4}(#:138,708)(126,708)(126,746){5}
wire [1:0] w12;    //: /sn:0 {0}(#:358,737)(358,768)(311,768){1}
//: {2}(309,766)(309,718)(376,718)(#:376,696){3}
//: {4}(309,770)(309,793)(330,793)(330,795){5}
wire w18;    //: /sn:0 {0}(673,594)(914,594){1}
//: {2}(918,594)(1344,594)(1344,572)(1357,572){3}
//: {4}(916,596)(916,649)(956,649)(956,618){5}
wire [1:0] w19;    //: /sn:0 {0}(#:295,1049)(295,979)(277,979)(277,942){1}
//: {2}(279,940)(344,940)(344,925){3}
//: {4}(#:277,938)(277,877)(330,877)(#:330,816){5}
wire w63;    //: /sn:0 {0}(382,418)(376,418)(376,416)(369,416){1}
//: {2}(367,414)(367,385)(1041,385){3}
//: {4}(365,416)(363,416)(363,412)(118,412){5}
//: {6}(116,410)(116,374)(204,374)(204,352)(166,352){7}
//: {8}(164,350)(164,232)(89,232)(89,195)(99,195){9}
//: {10}(162,352)(160,352){11}
//: {12}(116,414)(116,607)(108,607)(108,803){13}
//: {14}(110,805)(223,805){15}
//: {16}(227,805)(293,805){17}
//: {18}(225,807)(225,853)(479,853){19}
//: {20}(481,851)(481,806){21}
//: {22}(483,804)(490,804){23}
//: {24}(481,802)(481,745)(685,745)(685,735){25}
//: {26}(687,733)(705,733){27}
//: {28}(685,731)(685,667)(829,667){29}
//: {30}(833,667)(1793,667){31}
//: {32}(831,665)(831,533)(895,533){33}
//: {34}(683,733)(678,733){35}
//: {36}(481,855)(481,921)(614,921){37}
//: {38}(106,805)(81,805){39}
//: {40}(79,803)(79,756)(89,756){41}
//: {42}(79,807)(79,842)(-2,842){43}
//: {44}(-4,840)(-4,819)(-368,819)(-368,734)(-358,734){45}
//: {46}(-6,842)(-16,842)(-16,857)(-4,857){47}
//: {48}(108,807)(108,1072){49}
//: {50}(110,1074)(188,1074)(188,1076)(254,1076){51}
//: {52}(108,1076)(108,1244){53}
//: {54}(110,1246)(290,1246){55}
//: {56}(294,1246)(465,1246)(465,1225)(468,1225){57}
//: {58}(292,1244)(292,1230)(296,1230){59}
//: {60}(108,1248)(108,1467)(346,1467){61}
wire [1:0] w23;    //: /sn:0 {0}(#:823,136)(823,121){1}
wire [1:0] w10;    //: /sn:0 {0}(#:126,767)(126,782)(-55,782)(-55,930){1}
//: {2}(#:-53,932)(-32,932)(-32,917){3}
//: {4}(-55,934)(-55,1418)(506,1418)(506,1369)(#:498,1369){5}
wire [1:0] w24;    //: /sn:0 {0}(#:721,136)(721,121){1}
wire [1:0] w21;    //: /sn:0 {0}(#:506,1049)(506,1040)(524,1040)(524,944){1}
//: {2}(526,942)(527,942)(#:527,815){3}
//: {4}(522,942)(444,942)(444,925){5}
wire w31;    //: /sn:0 {0}(422,1472)(850,1472)(850,406){1}
//: {2}(852,404)(867,404)(867,374){3}
//: {4}(850,402)(850,293){5}
//: {6}(850,289)(850,268)(847,268)(847,257){7}
//: {8}(848,291)(836,291)(836,-96)(124,-96)(124,25)(141,25){9}
wire w1;    //: /sn:0 {0}(217,294)(248,294)(248,297)(258,297){1}
//: {2}(262,297)(281,297)(281,298)(300,298){3}
//: {4}(260,295)(260,192)(656,192){5}
wire [7:0] w32;    //: /sn:0 {0}(#:557,696)(557,750)(681,750)(681,765){1}
wire w53;    //: /sn:0 {0}(932,544)(932,562)(982,562)(982,574)(1122,574){1}
//: {2}(1126,574)(1243,574)(1243,381){3}
//: {4}(1243,377)(1243,373)(1371,373)(1371,385){5}
//: {6}(1241,379)(1165,379)(1165,390)(1117,390){7}
//: {8}(1124,572)(1124,535){9}
wire w46;    //: /sn:0 {0}(49,1172)(122,1172)(122,1139)(133,1139){1}
wire w17;    //: /sn:0 {0}(673,574)(858,574)(858,562)(917,562)(917,513)(932,513)(932,523){1}
wire [15:0] w27;    //: /sn:0 {0}(#:675,1066)(689,1066)(689,1073)(785,1073)(785,1554)(456,1554){1}
//: {2}(454,1552)(#:454,1531){3}
//: {4}(452,1554)(#:383,1554)(#:383,1478){5}
wire w44;    //: /sn:0 {0}(761,993)(905,993)(905,1572)(-308,1572)(-308,791)(-302,791)(-302,779)(-321,779)(-321,745){1}
wire [15:0] w28;    //: /sn:0 {0}(#:497,1146)(497,1169)(505,1169)(505,1190){1}
//: {2}(#:507,1192)(712,1192)(712,1176){3}
//: {4}(505,1194)(505,1215){5}
wire [15:0] w33;    //: /sn:0 {0}(#:333,1220)(333,1198){1}
//: {2}(333,1194)(333,1174){3}
//: {4}(335,1172)(639,1172)(639,1183)(1255,1183)(1255,412)(#:1270,412){5}
//: {6}(333,1170)(333,1159)(325,1159)(#:325,1146){7}
//: {8}(#:331,1196)(227,1196)(227,1178){9}
wire w35;    //: /sn:0 {0}(287,48)(287,65)(276,65)(276,4){1}
//: {2}(278,2)(309,2)(309,33)(1946,33)(1946,713)(1826,713)(1826,723){3}
//: {4}(1828,725)(1830,725)(1830,678){5}
//: {6}(1824,725)(1681,725)(1681,713)(1618,713)(1618,696){7}
//: {8}(274,2)(233,2){9}
//: {10}(231,0)(231,-32)(131,-32)(131,20)(141,20){11}
//: {12}(231,4)(231,25){13}
wire [7:0] w14;    //: /sn:0 {0}(#:637,869)(637,810)(691,810)(#:691,794){1}
wire w45;    //: /sn:0 {0}(740,990)(661,990){1}
//: {2}(657,990)(647,990)(647,1005)(678,1005)(678,1599)(77,1599)(77,1289)(196,1289){3}
//: {4}(659,992)(659,1033){5}
wire w49;    //: /sn:0 {0}(1078,396)(1078,411)(1141,411){1}
//: {2}(1145,411)(1162,411)(1162,397){3}
//: {4}(1143,413)(1143,588)(1357,588){5}
wire [15:0] w41;    //: /sn:0 {0}(#:642,875)(642,896)(651,896)(651,911){1}
wire [7:0] w2;    //: /sn:0 {0}(#:493,105)(493,63)(625,63){1}
//: {2}(629,63)(1956,63){3}
//: {4}(627,61)(627,2){5}
wire w48;    //: /sn:0 {0}(544,1230)(562,1230)(562,1281){1}
//: {2}(564,1283)(803,1283)(803,407)(809,407){3}
//: {4}(813,407)(827,407)(827,376){5}
//: {6}(811,405)(811,272)(800,272)(800,257){7}
//: {8}(560,1283)(377,1283)(377,1235)(372,1235){9}
wire [15:0] w47;    //: /sn:0 {0}(#:333,1241)(#:333,1255)(209,1255)(209,1273){1}
wire [7:0] w15;    //: /sn:0 {0}(#:612,696)(612,711){1}
wire w61;    //: /sn:0 {0}(908,175)(923,175){1}
wire w38;    //: /sn:0 {0}(1869,662)(1891,662)(1891,335)(1139,335)(1139,380)(1129,380){1}
//: {2}(1127,378)(1127,356)(969,356){3}
//: {4}(965,356)(480,356)(480,409){5}
//: {6}(482,411)(579,411)(579,327){7}
//: {8}(581,325)(1012,325)(1012,684){9}
//: {10}(1010,686)(1008,686)(1008,716)(789,716)(789,728)(781,728){11}
//: {12}(1012,688)(1012,799)(895,799){13}
//: {14}(891,799)(586,799){15}
//: {16}(582,799)(566,799){17}
//: {18}(584,801)(584,821){19}
//: {20}(582,823)(381,823)(381,802){21}
//: {22}(381,798)(381,751)(223,751){23}
//: {24}(219,751)(179,751){25}
//: {26}(177,749)(177,729)(-282,729){27}
//: {28}(175,751)(165,751){29}
//: {30}(221,753)(221,852)(72,852){31}
//: {32}(379,800)(369,800){33}
//: {34}(584,825)(584,1182)(595,1182)(595,1201){35}
//: {36}(597,1203)(598,1203)(598,1462)(422,1462){37}
//: {38}(593,1203)(555,1203){39}
//: {40}(551,1203)(376,1203)(376,1225)(372,1225){41}
//: {42}(553,1205)(553,1220)(544,1220){43}
//: {44}(893,801)(893,916)(690,916){45}
//: {46}(50:579,323)(579,306){47}
//: {48}(478,411)(474,411)(474,413)(458,413){49}
//: {50}(967,358)(967,517)(981,517)(981,528)(971,528){51}
//: {52}(1125,380)(1117,380){53}
wire w55;    //: /sn:0 {0}(1843,522)(1843,587)(1830,587)(1830,595){1}
//: {2}(1828,597)(1818,597)(1818,572)(1740,572){3}
//: {4}(1830,599)(1830,657){5}
wire w43;    //: /sn:0 {0}(221,54)(221,97)(276,97)(276,105){1}
wire [15:0] w26;    //: /sn:0 {0}(#:219,1302)(219,1316)(316,1316){1}
//: {2}(320,1316)(368,1316)(#:368,1331){3}
//: {4}(318,1318)(318,1345)(201,1345)(201,1361)(186,1361)(#:186,1349){5}
wire w9;    //: /sn:0 {0}(370,516)(370,493){1}
//: {2}(372,491)(388,491)(388,489)(410,489){3}
//: {4}(368,491)(51,491)(51,781)(668,781){5}
wire w40;    //: /sn:0 {0}(259,725)(259,738)(284,738){1}
//: {2}(286,736)(286,714)(284,714)(284,696){3}
//: {4}(286,740)(286,796)(33,796)(33,847){5}
wire w51;    //: /sn:0 {0}(1464,433)(1474,433)(1474,402){1}
//: {2}(1476,400)(1486,400)(1486,394)(1525,394)(1525,405)(1552,405)(1552,398){3}
//: {4}(1474,398)(1474,364)(1078,364)(1078,375){5}
//: enddecls

  //: GROUND g164 (w59) @(164,5) /sn:0 /w:[ 1 ]
  //: DIP g116 (w11) @(328,1275) /sn:0 /w:[ 0 ] /st:0 /dn:1
  _GGCLOCK_P200_0_50 g8 (.Z(w63));   //: @(147,352) /sn:0 /w:[ 11 ] /omega:200 /phi:0 /duty:50
  Instruction_Fetch g4 (.PC_in(w4), .EN(w1), .IR_OUT(w22));   //: @(301, 273) /sz:(200, 56) /sn:0 /p:[ Ti0>0 Li0>3 Bo0<0 ]
  //: joint g157 (w54) @(190, 192) /w:[ 2 4 6 1 ]
  //: joint g17 (w63) @(116, 412) /w:[ 5 6 -1 12 ]
  //: LED g137 (w53) @(1124,528) /sn:0 /w:[ 9 ] /type:0
  //: LED g30 (w22) @(532,347) /sn:0 /w:[ 3 ] /type:1
  //: LED g74 (w36) @(224,1399) /sn:0 /w:[ 5 ] /type:3
  //: joint g92 (w38) @(221, 751) /w:[ 23 -1 24 30 ]
  //: joint g1 (w63) @(164, 352) /w:[ 7 8 10 -1 ]
  jump_module g130 (.JNE_enable(w18), .Status_flag(w49), .offset_enable(w55));   //: @(1358, 556) /sz:(381, 80) /sn:0 /p:[ Li0>3 Li1>5 Ro0<3 ]
  //: LED g77 (w48) @(827,369) /sn:0 /w:[ 5 ] /type:0
  //: LED g111 (w16) @(193,1093) /sn:0 /w:[ 9 ] /type:0
  //: joint g144 (w55) @(1830, 597) /w:[ -1 1 2 4 ]
  _GGREG16 #(10, 10, 20) g51 (.Q(w47), .D(w33), .EN(~w48), .CLR(w38), .CK(w63));   //: @(333,1230) /sn:0 /w:[ 0 0 9 41 59 ]
  _GGAND2 #(6) g161 (.I0(w35), .I1(w31), .Z(w60));   //: @(152,23) /sn:0 /w:[ 11 9 0 ]
  _GGREG #(10, 10, 20) g70 (.Q(w56), .D(w29), .EN(~w30), .CLR(w38), .CK(w63));   //: @(742,733) /sn:0 /w:[ 3 5 13 11 27 ]
  //: joint g10 (w7) @(687, 404) /w:[ 4 6 -1 3 ]
  //: LED g149 (w55) @(1843,515) /sn:0 /w:[ 0 ] /type:0
  //: joint g25 (w30) @(125, 615) /w:[ 28 27 -1 30 ]
  //: LED g65 (w34) @(686,1285) /sn:0 /w:[ 3 ] /type:3
  //: joint g103 (w27) @(454, 1554) /w:[ 1 2 4 -1 ]
  //: joint g64 (w28) @(505, 1192) /w:[ 2 1 -1 4 ]
  //: joint g49 (w63) @(108, 1074) /w:[ 50 49 -1 52 ]
  //: LED g72 (w40) @(259,718) /sn:0 /w:[ 0 ] /type:0
  //: joint g142 (w18) @(916, 594) /w:[ 2 -1 1 4 ]
  //: LED g136 (w49) @(1162,390) /sn:0 /w:[ 3 ] /type:0
  Instruction_Decode g6 (.IR_IN(w6), .EN(w30), .IN2_User(w9), .ALU_MODE(w37), .ALU_EN(w40), .Reg1(w12), .Reg2(w13), .Imm2(w32), .MemAddr2(w15), .RW1(w29), .Cmp_EN(w17), .Jmp_EN(w18), .RR(w20), .HLT(w58));   //: @(209, 517) /sz:(463, 178) /sn:0 /p:[ Li0>5 Li1>31 To0<0 Bo0<0 Bo1<3 Bo2<3 Bo3<3 Bo4<0 Bo5<0 Ro0<0 Ro1<0 Ro2<0 Ro3<0 Ro4<0 ]
  //: joint g124 (w63) @(-4, 842) /w:[ 43 44 46 -1 ]
  //: joint g35 (w12) @(309, 768) /w:[ 1 2 -1 4 ]
  //: joint g7 (w6) @(407, 479) /w:[ 2 1 4 -1 ]
  //: joint g56 (w63) @(292, 1246) /w:[ 56 58 55 -1 ]
  //: LED g58 (w27) @(454,1524) /sn:0 /w:[ 3 ] /type:3
  //: joint g98 (w56) @(61, 1106) /w:[ -1 6 5 8 ]
  //: LED g67 (w26) @(186,1342) /sn:0 /w:[ 5 ] /type:3
  //: joint g85 (w30) @(756, 757) /w:[ 8 14 -1 7 ]
  //: joint g126 (w16) @(218, 1119) /w:[ 4 6 -1 3 ]
  //: joint g33 (w30) @(756, 405) /w:[ 20 -1 22 19 ]
  //: joint g54 (w38) @(553, 1203) /w:[ 39 -1 40 42 ]
  Register_File g40 (.Addr2(w21), .Write_Data(w25), .Addr1(w19), .RW1(w16), .CLK(w63), .CLR(w0), .Data_out2(w28), .Data_out1(w33));   //: @(255, 1050) /sz:(291, 95) /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>0 Li0>5 Li1>51 Ri0>15 Bo0<0 Bo1<7 ]
  _GGREG16 #(10, 10, 20) g52 (.Q(w34), .D(w28), .EN(~w48), .CLR(w38), .CK(w63));   //: @(505,1225) /sn:0 /w:[ 5 5 0 43 57 ]
  //: joint g81 (w38) @(584, 823) /w:[ -1 19 20 34 ]
  //: joint g163 (w35) @(276, 2) /w:[ 2 -1 8 1 ]
  //: DIP g132 (w52) @(1187,310) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: joint g12 (w0) @(388, 55) /w:[ 3 4 -1 10 ]
  //: joint g108 (w7) @(638, 422) /w:[ 2 -1 1 8 ]
  Comparator_16Bit g131 (.EN(w53), .Reg1(w33), .Reg2(w52), .Out(w51));   //: @(1271, 386) /sz:(192, 115) /sn:0 /p:[ Ti0>5 Li0>5 Li1>1 Ro0<0 ]
  //: LED g106 (w25) @(352,991) /sn:0 /w:[ 5 ] /type:3
  //: joint g96 (w10) @(-55, 932) /w:[ 2 1 -1 4 ]
  //: joint g19 (w48) @(811, 407) /w:[ 4 6 3 -1 ]
  //: joint g114 (w50) @(21, 1133) /w:[ 5 -1 6 12 ]
  //: joint g117 (w20) @(1055, 654) /w:[ 2 4 1 -1 ]
  //: joint g78 (w0) @(579, 201) /w:[ 1 2 -1 12 ]
  //: joint g125 (w42) @(689, 1006) /w:[ 7 -1 8 10 ]
  //: joint g155 (w35) @(1826, 725) /w:[ 4 3 6 -1 ]
  //: LED g63 (w28) @(712,1169) /sn:0 /w:[ 3 ] /type:3
  //: LED g93 (w50) @(65,927) /sn:0 /w:[ 0 ] /type:0
  //: joint g100 (w38) @(893, 799) /w:[ 13 -1 14 44 ]
  _GGMUX2x16 #(8, 8) g105 (.I0(w42), .I1(w27), .S(w45), .Z(w25));   //: @(659,1056) /sn:0 /R:3 /w:[ 11 0 5 3 ] /ss:0 /do:0
  _GGAND2 #(6) g113 (.I0(w50), .I1(w7), .Z(w46));   //: @(39,1172) /sn:0 /w:[ 13 9 0 ]
  Program_Counter g0 (.Offset_IN(w2), .CLR(w0), .Offset_EN(w43), .CLK(w54), .PC_OUT(w4));   //: @(213, 106) /sz:(357, 74) /sn:0 /p:[ Ti0>0 Ti1>11 Ti2>1 Li0>5 Bo0<5 ]
  //: joint g38 (w22) @(407, 381) /w:[ 2 1 -1 4 ]
  assign w41 = {w8, w14}; //: CONCAT g43  @(642,874) /sn:0 /R:3 /w:[ 0 1 0 ] /dr:0 /tp:0 /drp:1
  //: joint g101 (w30) @(756, 835) /w:[ -1 6 5 32 ]
  _GGREG16 #(10, 10, 20) g48 (.Q(w27), .D(w36), .EN(~w31), .CLR(w38), .CK(w63));   //: @(383,1467) /sn:0 /w:[ 5 0 0 37 61 ]
  //: joint g37 (w13) @(527, 751) /w:[ -1 2 1 4 ]
  //: joint g80 (w1) @(260, 297) /w:[ 2 4 1 -1 ]
  //: joint g122 (w38) @(177, 751) /w:[ 25 26 28 -1 ]
  _GGREG #(10, 10, 20) g120 (.Q(w44), .D(w20), .EN(~w30), .CLR(w38), .CK(w63));   //: @(-321,734) /sn:0 /w:[ 1 5 43 27 45 ]
  //: LED g95 (w10) @(-32,910) /sn:0 /w:[ 3 ] /type:1
  //: joint g76 (w26) @(318, 1316) /w:[ 2 -1 1 4 ]
  //: DIP g170 (w62) @(891,739) /sn:0 /w:[ 0 ] /st:7 /dn:1
  //: joint g152 (w38) @(967, 356) /w:[ 3 -1 4 50 ]
  //: joint g44 (w63) @(108, 805) /w:[ 14 13 38 48 ]
  //: joint g75 (w36) @(383, 1439) /w:[ -1 2 4 1 ]
  _GGAND2 #(6) g159 (.I0(~w58), .I1(w63), .Z(w54));   //: @(110,193) /sn:0 /w:[ 3 9 7 ]
  //: SWITCH g3 (w0) @(361,-64) /sn:0 /w:[ 7 ] /st:1 /dn:1
  //: LED g16 (w6) @(564,439) /sn:0 /w:[ 3 ] /type:1
  //: LED g47 (w39) @(488,1407) /sn:0 /R:2 /w:[ 0 ] /type:0
  _GGREG #(10, 10, 20) g143 (.Q(w35), .D(w55), .EN(~w30), .CLR(w38), .CK(w63));   //: @(1830,667) /sn:0 /w:[ 5 5 17 0 31 ]
  //: joint g26 (w63) @(225, 805) /w:[ 16 -1 15 18 ]
  //: joint g90 (w40) @(286, 738) /w:[ -1 2 1 4 ]
  _GGMUX2 #(8, 8) g109 (.I0(w46), .I1(w56), .S(w56), .Z(w16));   //: @(149,1129) /sn:0 /R:1 /w:[ 1 9 0 0 ] /ss:0 /do:0
  //: LED g158 (w35) @(287,41) /sn:0 /w:[ 0 ] /type:0
  //: LED g2 (w2) @(627,-5) /sn:0 /w:[ 5 ] /type:3
  //: joint g128 (w63) @(367, 416) /w:[ 1 2 4 -1 ]
  _GGREG2 #(10, 10, 20) g23 (.Q(w19), .D(w12), .EN(~w30), .CLR(w38), .CK(w63));   //: @(330,805) /sn:0 /w:[ 5 5 37 33 17 ]
  //: joint g91 (w63) @(79, 805) /w:[ 39 40 -1 42 ]
  _GGMUX2x16 #(8, 8) g104 (.I0(w47), .I1(w11), .S(w45), .Z(w26));   //: @(219,1289) /sn:0 /w:[ 1 1 3 0 ] /ss:0 /do:0
  //: LED g141 (w18) @(956,611) /sn:0 /w:[ 5 ] /type:0
  _GGREG2 #(10, 10, 20) g24 (.Q(w21), .D(w13), .EN(~w30), .CLR(w38), .CK(w63));   //: @(527,804) /sn:0 /w:[ 3 5 35 17 23 ]
  //: LED g39 (w30) @(151,591) /sn:0 /w:[ 29 ] /type:0
  //: joint g86 (w37) @(140, 708) /w:[ 1 2 4 -1 ]
  _GGREG #(10, 10, 20) g127 (.Q(w49), .D(w51), .EN(~w53), .CLR(w38), .CK(w63));   //: @(1078,385) /sn:0 /w:[ 0 5 7 53 3 ]
  //: joint g29 (w38) @(584, 799) /w:[ 15 -1 16 18 ]
  _GGREG16 #(10, 10, 20) g60 (.Q(w42), .D(w41), .EN(~w30), .CLR(w38), .CK(w63));   //: @(651,921) /sn:0 /w:[ 9 1 33 45 37 ]
  //: joint g110 (w56) @(-13, 1006) /w:[ 1 2 -1 4 ]
  //: joint g121 (w50) @(-11, 1296) /w:[ 8 7 -1 10 ]
  //: LED g168 (w58) @(42,307) /sn:0 /w:[ 5 ] /type:0
  //: LED g18 (w7) @(687,370) /sn:0 /w:[ 7 ] /type:0
  //: joint g82 (w29) @(742, 540) /w:[ -1 2 1 4 ]
  //: LED g119 (w20) @(1088,571) /sn:0 /w:[ 3 ] /type:0
  //: joint g94 (w50) @(33, 945) /w:[ 1 2 -1 4 ]
  //: SWITCH g173 (w54) @(217,232) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: joint g166 (w35) @(231, 2) /w:[ 9 10 -1 12 ]
  assign w2 = w42[7:0]; //: TAP g154 @(1959,63) /sn:0 /R:2 /w:[ 3 3 4 ] /ss:0
  //: joint g107 (w25) @(412, 1033) /w:[ -1 2 4 1 ]
  //: joint g172 (w9) @(370, 491) /w:[ 2 -1 4 1 ]
  //: joint g50 (w21) @(524, 942) /w:[ 2 -1 4 1 ]
  Control_Unit g9 (.OP1(w24), .OP2(w23), .CLK(w54), .EN_Decoder(w1), .CLR(w0), .EN1(w7), .EN2(w30), .EN3(w48), .EN4(w31), .OP_Forwarding(w61));   //: @(657, 137) /sz:(250, 119) /sn:0 /p:[ Ti0>0 Ti1>0 Li0>3 Li1>5 Li2>0 Bo0<5 Bo1<25 Bo2<7 Bo3<7 Ro0<0 ]
  //: joint g133 (w33) @(333, 1172) /w:[ 4 6 -1 3 ]
  //: LED g68 (w37) @(140,674) /sn:0 /w:[ 3 ] /type:1
  _GGREG #(10, 10, 20) g73 (.Q(w50), .D(w40), .EN(~w30), .CLR(w38), .CK(w63));   //: @(33,857) /sn:0 /w:[ 3 5 0 31 47 ]
  _GGMUX2x8 #(8, 8) g169 (.I0(w32), .I1(w62), .S(w9), .Z(w14));   //: @(691,781) /sn:0 /w:[ 1 1 5 1 ] /ss:0 /do:0
  //: joint g31 (w30) @(574, 835) /w:[ 4 34 3 -1 ]
  //: joint g22 (w38) @(579, 325) /w:[ 8 46 -1 7 ]
  //: LED g59 (w42) @(770,952) /sn:0 /w:[ 0 ] /type:3
  //: LED g71 (w29) @(742,518) /sn:0 /w:[ 3 ] /type:0
  //: joint g102 (w63) @(481, 853) /w:[ -1 20 19 36 ]
  //: joint g87 (w38) @(1012, 686) /w:[ -1 9 10 12 ]
  _GGAND2 #(6) g99 (.I0(w44), .I1(w16), .Z(w45));   //: @(750,990) /sn:0 /R:2 /w:[ 0 7 0 ]
  //: joint g83 (w63) @(481, 804) /w:[ 22 24 -1 21 ]
  //: joint g45 (w31) @(850, 404) /w:[ 2 4 -1 1 ]
  //: LED g36 (w13) @(417,734) /sn:0 /w:[ 0 ] /type:1
  //: joint g41 (w19) @(277, 940) /w:[ 2 4 -1 1 ]
  //: SWITCH g42 (w8) @(696,861) /sn:0 /R:2 /w:[ 0 ] /st:0 /dn:1
  _GGREG2 #(10, 10, 20) g69 (.Q(w10), .D(w37), .EN(~w30), .CLR(w38), .CK(w63));   //: @(126,756) /sn:0 /w:[ 0 5 41 29 41 ]
  //: joint g156 (w2) @(627, 63) /w:[ 2 4 1 -1 ]
  //: joint g138 (w53) @(1124, 574) /w:[ 2 8 1 -1 ]
  //: joint g167 (w58) @(73, 339) /w:[ 2 -1 4 1 ]
  //: joint g151 (w30) @(788, 745) /w:[ 10 12 -1 9 ]
  //: joint g66 (w34) @(472, 1305) /w:[ 2 4 -1 1 ]
  //: joint g153 (w42) @(770, 1003) /w:[ 2 1 -1 6 ]
  //: joint g146 (w30) @(756, 513) /w:[ 16 18 -1 15 ]
  //: joint g162 (w0) @(388, -9) /w:[ -1 6 8 5 ]
  //: LED g34 (w12) @(358,730) /sn:0 /w:[ 0 ] /type:1
  //: LED g28 (w21) @(444,918) /sn:0 /w:[ 5 ] /type:1
  ALU g46 (.IN2(w34), .IN1(w26), .EN(w50), .MODE(w10), .OF(w39), .OUT(w36));   //: @(349, 1332) /sz:(148, 53) /sn:0 /p:[ Ti0>0 Ti1>3 Li0>11 Ri0>5 Bo0<1 Bo1<3 ]
  //: joint g57 (w63) @(108, 1246) /w:[ 54 53 -1 60 ]
  //: joint g11 (w30) @(742, 405) /w:[ 23 24 -1 26 ]
  //: joint g150 (w63) @(831, 667) /w:[ 30 32 29 -1 ]
  //: joint g14 (w0) @(579, 217) /w:[ 14 13 -1 16 ]
  //: joint g84 (w63) @(685, 733) /w:[ 26 28 34 25 ]
  //: LED g118 (w50) @(34,1280) /sn:0 /w:[ 9 ] /type:0
  _GGNBUF #(2) g5 (.I(w0), .Z(w1));   //: @(207,294) /sn:0 /w:[ 9 0 ]
  //: joint g112 (w16) @(193, 1128) /w:[ 2 8 1 -1 ]
  //: joint g123 (w30) @(152, 776) /w:[ 40 42 39 -1 ]
  //: joint g21 (w4) @(391, 263) /w:[ 2 4 -1 1 ]
  //: LED g61 (w33) @(227,1171) /sn:0 /w:[ 9 ] /type:3
  //: LED g79 (w31) @(867,367) /sn:0 /w:[ 3 ] /type:0
  //: LED g20 (w4) @(432,241) /sn:0 /w:[ 3 ] /type:3
  //: LED g32 (w30) @(776,371) /sn:0 /w:[ 21 ] /type:0
  //: joint g115 (w45) @(659, 990) /w:[ 1 -1 2 4 ]
  //: LED g97 (w56) @(81,1103) /sn:0 /R:2 /w:[ 7 ] /type:0
  //: LED g134 (w51) @(1552,391) /sn:0 /w:[ 3 ] /type:0
  //: joint g145 (w38) @(1127, 380) /w:[ 1 2 52 -1 ]
  _GGREG #(10, 10, 20) g148 (.Q(w53), .D(w17), .EN(~w30), .CLR(w38), .CK(w63));   //: @(932,533) /sn:0 /w:[ 0 1 11 51 33 ]
  //: joint g89 (w30) @(377, 835) /w:[ 2 36 38 1 ]
  _GGREG16 #(10, 10, 20) g15 (.Q(w6), .D(w22), .EN(~w7), .CLR(w38), .CK(w63));   //: @(419,418) /sn:0 /w:[ 0 5 0 49 0 ]
  //: joint g129 (w38) @(480, 411) /w:[ 6 5 48 -1 ]
  //: LED g27 (w19) @(344,918) /sn:0 /w:[ 3 ] /type:1
  //: LED g147 (w35) @(1618,689) /sn:0 /w:[ 7 ] /type:0
  //: joint g165 (w31) @(850, 291) /w:[ -1 6 8 5 ]
  //: LED g171 (w9) @(417,489) /sn:0 /R:3 /w:[ 3 ] /type:0
  //: joint g62 (w33) @(333, 1196) /w:[ -1 2 8 1 ]
  _GGMUX2 #(8, 8) g160 (.I0(w59), .I1(w35), .S(w60), .Z(w43));   //: @(221,41) /sn:0 /w:[ 0 13 1 0 ] /ss:0 /do:0
  //: joint g88 (w38) @(381, 800) /w:[ -1 22 32 21 ]
  //: joint g55 (w38) @(595, 1203) /w:[ 36 35 38 -1 ]
  //: joint g53 (w48) @(562, 1283) /w:[ 2 1 8 -1 ]
  _GGNBUF #(2) g13 (.I(w0), .Z(w38));   //: @(579,296) /sn:0 /R:3 /w:[ 17 47 ]
  //: joint g135 (w51) @(1474, 400) /w:[ 2 4 -1 1 ]
  //: joint g140 (w49) @(1143, 411) /w:[ 2 -1 1 4 ]
  //: joint g139 (w53) @(1243, 379) /w:[ -1 4 6 3 ]

endmodule
//: /netlistEnd

//: /netlistBegin Comparator_2bit
module Comparator_2bit(Reg2, Out, Reg1);
//: interface  /sz:(133, 95) /bd:[ Ti0>Reg2[1:0](105/133) Ti1>Reg1[1:0](18/133) Bo0<Out(62/133) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
output Out;    //: /sn:0 {0}(382,428)(382,467)(396,467){1}
input [1:0] Reg1;    //: /sn:0 {0}(#:462,105)(462,154)(423,154){1}
//: {2}(422,154)(349,154){3}
//: {4}(348,154)(#:246,154){5}
input [1:0] Reg2;    //: /sn:0 {0}(#:490,139)(490,218)(427,218){1}
//: {2}(426,218)(357,218){3}
//: {4}(356,218)(#:249,218){5}
wire w4;    //: /sn:0 {0}(423,158)(423,166)(421,166)(421,303){1}
wire w3;    //: /sn:0 {0}(427,222)(427,230)(426,230)(426,303){1}
wire w0;    //: /sn:0 {0}(357,222)(357,232)(354,232)(354,301){1}
wire w1;    //: /sn:0 {0}(349,158)(349,301){1}
wire w2;    //: /sn:0 {0}(380,407)(380,333)(351,333)(351,322){1}
wire w5;    //: /sn:0 {0}(385,407)(385,335)(423,335)(423,324){1}
//: enddecls

  _GGAND2 #(6) g8 (.I0(w5), .I1(w2), .Z(Out));   //: @(382,418) /sn:0 /R:3 /w:[ 0 0 0 ]
  assign w1 = Reg1[0]; //: TAP g4 @(349,152) /sn:0 /R:1 /w:[ 0 4 3 ] /ss:1
  _GGNXOR2 #(6) g3 (.I0(w3), .I1(w4), .Z(w5));   //: @(423,314) /sn:0 /R:3 /w:[ 1 1 1 ]
  _GGNXOR2 #(6) g2 (.I0(w0), .I1(w1), .Z(w2));   //: @(351,312) /sn:0 /R:3 /w:[ 1 1 1 ]
  //: IN g1 (Reg2) @(247,218) /sn:0 /w:[ 5 ]
  //: LED g10 (Reg1) @(462,98) /sn:0 /w:[ 0 ] /type:1
  assign w4 = Reg1[1]; //: TAP g6 @(423,152) /sn:0 /R:1 /w:[ 0 2 1 ] /ss:1
  //: OUT g9 (Out) @(393,467) /sn:0 /w:[ 1 ]
  assign w3 = Reg2[1]; //: TAP g7 @(427,216) /sn:0 /R:1 /w:[ 0 2 1 ] /ss:1
  //: LED g11 (Reg2) @(490,132) /sn:0 /w:[ 0 ] /type:1
  assign w0 = Reg2[0]; //: TAP g5 @(357,216) /sn:0 /R:1 /w:[ 0 4 3 ] /ss:1
  //: IN g0 (Reg1) @(244,154) /sn:0 /w:[ 5 ]

endmodule
//: /netlistEnd

//: /netlistBegin Program_Counter
module Program_Counter(PC_OUT, Offset_IN, CLK, Offset_EN, CLR);
//: interface  /sz:(357, 74) /bd:[ Ti0>Offset_IN[7:0](280/357) Ti1>CLR(176/357) Ti2>Offset_EN(63/357) Li0>CLK(36/74) Bo0<PC_OUT[7:0](179/357) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
output [7:0] PC_OUT;    //: {0}(#:-1:427,387)(427,400)(#:494,400){1}
//: {2}(498,400)(551,400){3}
//: {4}(555,400)(692,400)(#:692,414){5}
//: {6}(553,398)(553,359){7}
//: {8}(496,398)(#:496,281){9}
input Offset_EN;    //: /sn:0 {0}(440,462)(450,462)(450,445)(332,445){1}
input [7:0] Offset_IN;    //: /sn:0 {0}(#:204,491)(204,528)(297,528){1}
//: {2}(301,528)(#:377,528){3}
//: {4}(299,526)(299,461){5}
supply0 w3;    //: /sn:0 {0}(535,275)(571,275)(571,294){1}
reg w1;    //: /sn:0 {0}(732,428)(776,428){1}
input CLR;    //: /sn:0 {0}(568,165)(568,205){1}
input CLK;    //: /sn:0 {0}(459,270)(377,270)(377,278){1}
reg [7:0] w5;    //: /sn:0 {0}(#:725,346)(725,404)(724,404)(724,414){1}
wire [7:0] w7;    //: /sn:0 {0}(#:309,432)(309,393)(310,393)(310,360){1}
//: {2}(310,356)(310,234)(496,234)(#:496,260){3}
//: {4}(#:308,358)(250,358)(250,319){5}
wire [7:0] w8;    //: /sn:0 {0}(#:319,461)(319,508)(708,508)(#:708,443){1}
wire w2;    //: /sn:0 {0}(568,221)(568,253){1}
//: {2}(570,255)(592,255)(592,234){3}
//: {4}(568,257)(568,265)(535,265){5}
wire w9;    //: /sn:0 {0}(613,428)(684,428){1}
//: enddecls

  //: LED g4 (w9) @(606,428) /sn:0 /R:1 /w:[ 0 ] /type:0
  //: OUT g8 (PC_OUT) @(427,390) /sn:0 /R:1 /w:[ 0 ]
  //: SWITCH g3 (w1) @(794,428) /sn:0 /R:2 /w:[ 1 ] /st:0 /dn:1
  //: LED g16 (w7) @(250,312) /sn:0 /w:[ 5 ] /type:3
  //: joint g17 (w7) @(310, 358) /w:[ -1 2 4 1 ]
  //: joint g2 (PC_OUT) @(496, 400) /w:[ 2 8 1 -1 ]
  _GGADD8 #(68, 70, 62, 64) g1 (.A(PC_OUT), .B(w5), .S(w8), .CI(w1), .CO(w9));   //: @(708,430) /sn:0 /w:[ 5 1 1 0 1 ]
  //: LED g18 (PC_OUT) @(553,352) /sn:0 /w:[ 7 ] /type:3
  _GGMUX2x8 #(8, 8) g10 (.I0(w8), .I1(Offset_IN), .S(Offset_EN), .Z(w7));   //: @(309,445) /sn:0 /R:2 /w:[ 0 5 1 0 ] /ss:0 /do:0
  //: IN g6 (Offset_IN) @(379,528) /sn:0 /R:2 /w:[ 3 ]
  //: GROUND g9 (w3) @(571,300) /sn:0 /w:[ 1 ]
  //: IN g7 (CLK) @(377,280) /sn:0 /R:1 /w:[ 1 ]
  //: IN g12 (Offset_EN) @(438,462) /sn:0 /w:[ 0 ]
  //: DIP g5 (w5) @(725,336) /sn:0 /w:[ 0 ] /st:1 /dn:1
  //: IN g11 (CLR) @(568,163) /sn:0 /R:3 /w:[ 0 ]
  //: LED g14 (w2) @(592,227) /sn:0 /w:[ 3 ] /type:0
  //: joint g19 (PC_OUT) @(553, 400) /w:[ 4 6 3 -1 ]
  //: joint g21 (Offset_IN) @(299, 528) /w:[ 2 4 1 -1 ]
  //: LED g20 (Offset_IN) @(204,484) /sn:0 /w:[ 0 ] /type:3
  _GGREG8 #(10, 10, 20) g0 (.Q(PC_OUT), .D(w7), .EN(w3), .CLR(w2), .CK(CLK));   //: @(496,270) /sn:0 /w:[ 9 3 0 5 0 ]
  //: joint g15 (w2) @(568, 255) /w:[ 2 1 -1 4 ]
  _GGNBUF #(2) g13 (.I(CLR), .Z(w2));   //: @(568,211) /sn:0 /R:3 /w:[ 1 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin Comparator_16Bit
module Comparator_16Bit(Reg2, EN, Out, Reg1);
//: interface  /sz:(192, 115) /bd:[ Ti0>EN(100/192) Li0>Reg1[15:0](26/115) Li1>Reg2[15:0](83/115) Ro0<Out(47/115) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
output Out;    //: /sn:0 {0}(665,375)(665,418)(685,418){1}
input [15:0] Reg1;    //: /sn:0 {0}(#:62,-9)(105,-9){1}
input EN;    //: /sn:0 {0}(-10,-81)(20,-81){1}
//: {2}(24,-81)(113,-81)(113,-14){3}
//: {4}(22,-83)(22,-122)(-38,-122)(-38,-53)(12,-53)(12,21)(85,21)(85,52){5}
input [15:0] Reg2;    //: /sn:0 {0}(77,57)(38,57)(38,58)(#:11,58){1}
wire w6;    //: /sn:0 {0}(642,354)(642,309)(421,309)(421,165){1}
wire w13;    //: /sn:0 {0}(647,354)(647,303)(528,303)(528,161){1}
wire w16;    //: /sn:0 {0}(600,-4)(600,4)(598,4)(598,142){1}
wire w7;    //: /sn:0 {0}(347,160)(347,316)(637,316)(637,354){1}
wire w58;    //: /sn:0 {0}(702,354)(702,342)(1510,342)(1510,167){1}
wire w34;    //: /sn:0 {0}(1152,-4)(1152,4)(1150,4)(1150,147){1}
wire w50;    //: /sn:0 {0}(1256,-6)(1256,143){1}
wire w59;    //: /sn:0 {0}(1438,165)(1438,335)(697,335)(697,354){1}
wire w4;    //: /sn:0 {0}(239,-5)(239,3)(237,3)(237,140){1}
wire w25;    //: /sn:0 {0}(900,165)(900,303)(667,303)(667,354){1}
wire w62;    //: /sn:0 {0}(1436,-5)(1436,144){1}
wire [15:0] w39;    //: /sn:0 {0}(#:121,-9)(164,-9){1}
//: {2}(165,-9)(238,-9){3}
//: {4}(239,-9)(316,-9)(#:316,-8)(344,-8){5}
//: {6}(345,-8)(421,-8){7}
//: {8}(422,-8)(525,-8){9}
//: {10}(526,-8)(599,-8){11}
//: {12}(600,-8)(708,-8){13}
//: {14}(709,-8)(782,-8){15}
//: {16}(783,-8)(903,-8){17}
//: {18}(904,-8)(970,-8){19}
//: {20}(971,-8)(1078,-8){21}
//: {22}(1079,-8)(1151,-8){23}
//: {24}(1152,-8)(1227,-8)(#:1227,-10)(1255,-10){25}
//: {26}(1256,-10)(1329,-10){27}
//: {28}(1330,-10)(1407,-10)(#:1407,-9)(1435,-9){29}
//: {30}(1436,-9)(1509,-9){31}
//: {32}(1510,-9)(1609,-9)(#:1609,-28){33}
wire w56;    //: /sn:0 {0}(1444,65)(1444,75)(1441,75)(1441,144){1}
wire w3;    //: /sn:0 {0}(243,59)(243,67)(242,67)(242,140){1}
wire w0;    //: /sn:0 {0}(173,59)(173,69)(170,69)(170,138){1}
wire w22;    //: /sn:0 {0}(783,-4)(783,4)(778,4)(778,143){1}
wire w36;    //: /sn:0 {0}(692,354)(692,327)(1330,327)(1330,166){1}
wire w20;    //: /sn:0 {0}(780,164)(780,300)(662,300)(662,354){1}
wire w29;    //: /sn:0 {0}(1156,66)(1156,74)(1155,74)(1155,147){1}
wire w30;    //: /sn:0 {0}(1086,66)(1086,139)(1083,139)(1083,145){1}
wire w37;    //: /sn:0 {0}(687,354)(687,322)(1258,322)(1258,164){1}
wire w12;    //: /sn:0 {0}(652,354)(652,297)(600,297)(600,163){1}
wire w18;    //: /sn:0 {0}(714,62)(714,72)(711,72)(711,141){1}
wire w19;    //: /sn:0 {0}(534,61)(534,71)(531,71)(531,140){1}
wire w10;    //: /sn:0 {0}(422,-4)(422,4)(419,4)(419,144){1}
wire w23;    //: /sn:0 {0}(709,-4)(709,67)(706,67)(706,141){1}
wire w54;    //: /sn:0 {0}(1514,65)(1514,73)(1513,73)(1513,146){1}
wire w21;    //: /sn:0 {0}(657,354)(657,295)(708,295)(708,162){1}
wire w24;    //: /sn:0 {0}(672,354)(672,306)(972,306)(972,167){1}
wire w1;    //: /sn:0 {0}(165,-5)(165,138){1}
wire w31;    //: /sn:0 {0}(906,65)(906,75)(903,75)(903,144){1}
wire w32;    //: /sn:0 {0}(1152,168)(1152,317)(682,317)(682,354){1}
wire w53;    //: /sn:0 {0}(1330,-6)(1330,2)(1328,2)(1328,145){1}
wire w8;    //: /sn:0 {0}(345,-4)(345,139){1}
wire w52;    //: /sn:0 {0}(1334,64)(1334,72)(1333,72)(1333,145){1}
wire w17;    //: /sn:0 {0}(784,62)(784,70)(783,70)(783,143){1}
wire w27;    //: /sn:0 {0}(976,65)(976,73)(975,73)(975,146){1}
wire w28;    //: /sn:0 {0}(971,-4)(971,4)(970,4)(970,146){1}
wire w33;    //: /sn:0 {0}(677,354)(677,311)(1080,311)(1080,166){1}
wire w35;    //: /sn:0 {0}(1079,-4)(1079,42)(1078,42)(1078,145){1}
wire w14;    //: /sn:0 {0}(526,-4)(526,140){1}
wire w2;    //: /sn:0 {0}(627,354)(627,330)(167,330)(167,159){1}
wire w11;    //: /sn:0 {0}(353,60)(353,70)(350,70)(350,139){1}
wire w15;    //: /sn:0 {0}(604,61)(604,69)(603,69)(603,142){1}
wire w5;    //: /sn:0 {0}(239,161)(239,323)(632,323)(632,354){1}
wire w61;    //: /sn:0 {0}(1510,-5)(1510,3)(1508,3)(1508,146){1}
wire [15:0] w38;    //: /sn:0 {0}(#:93,57)(109,57)(109,55)(172,55){1}
//: {2}(173,55)(242,55){3}
//: {4}(243,55)(315,55)(#:315,56)(352,56){5}
//: {6}(353,56)(389,56)(389,59)(424,59){7}
//: {8}(425,59)(496,59)(#:496,57)(533,57){9}
//: {10}(534,57)(603,57){11}
//: {12}(604,57)(676,57)(#:676,58)(713,58){13}
//: {14}(714,58)(783,58){15}
//: {16}(784,58)(868,58)(#:868,61)(905,61){17}
//: {18}(906,61)(975,61){19}
//: {20}(976,61)(1048,61)(#:1048,62)(1085,62){21}
//: {22}(1086,62)(1155,62){23}
//: {24}(1156,62)(1184,62)(1184,60)(1263,60){25}
//: {26}(1264,60)(1333,60){27}
//: {28}(1334,60)(1413,60)(1413,61)(1443,61){29}
//: {30}(1444,61)(1513,61){31}
//: {32}(1514,61)(1651,61)(#:1651,28){33}
wire w9;    //: /sn:0 {0}(425,63)(425,71)(424,71)(424,144){1}
wire w26;    //: /sn:0 {0}(904,-4)(904,67)(898,67)(898,144){1}
wire w57;    //: /sn:0 {0}(1264,64)(1264,74)(1261,74)(1261,143){1}
//: enddecls

  assign w1 = w39[0]; //: TAP g4 @(165,-11) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  assign w27 = w38[9]; //: TAP g44 @(976,59) /sn:0 /R:1 /w:[ 0 19 20 ] /ss:1
  _GGAND16 #(34) g8 (.I0(w58), .I1(w59), .I2(w36), .I3(w37), .I4(w32), .I5(w33), .I6(w24), .I7(w25), .I8(w20), .I9(w21), .I10(w12), .I11(w13), .I12(w6), .I13(w7), .I14(w5), .I15(w2), .Z(Out));   //: @(665,365) /sn:0 /R:3 /w:[ 0 1 0 0 1 0 0 1 1 0 0 0 0 1 1 0 0 ]
  _GGNXOR2 #(6) g3 (.I0(w3), .I1(w4), .Z(w5));   //: @(239,151) /sn:0 /R:3 /w:[ 1 1 0 ]
  assign w9 = w38[3]; //: TAP g16 @(425,57) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  assign w35 = w39[10]; //: TAP g47 @(1079,-10) /sn:0 /R:1 /w:[ 0 21 22 ] /ss:1
  assign w11 = w38[2]; //: TAP g17 @(353,54) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  //: joint g26 (EN) @(22, -81) /w:[ 2 4 1 -1 ]
  _GGNXOR2 #(6) g2 (.I0(w0), .I1(w1), .Z(w2));   //: @(167,149) /sn:0 /R:3 /w:[ 1 1 1 ]
  _GGNXOR2 #(6) g23 (.I0(w19), .I1(w14), .Z(w13));   //: @(528,151) /sn:0 /R:3 /w:[ 1 1 1 ]
  assign w23 = w39[6]; //: TAP g30 @(709,-10) /sn:0 /R:1 /w:[ 0 13 14 ] /ss:1
  //: IN g1 (Reg2) @(9,58) /sn:0 /w:[ 1 ]
  _GGNXOR2 #(6) g39 (.I0(w31), .I1(w26), .Z(w25));   //: @(900,155) /sn:0 /R:3 /w:[ 1 1 0 ]
  assign w19 = w38[4]; //: TAP g29 @(534,55) /sn:0 /R:1 /w:[ 0 9 10 ] /ss:1
  assign w52 = w38[13]; //: TAP g60 @(1334,58) /sn:0 /R:1 /w:[ 0 27 28 ] /ss:1
  assign w16 = w39[5]; //: TAP g25 @(600,-10) /sn:0 /R:1 /w:[ 0 11 12 ] /ss:1
  _GGBUFIF16 #(4, 6) g10 (.Z(w39), .I(Reg1), .E(EN));   //: @(111,-9) /sn:0 /w:[ 0 1 3 ]
  assign w61 = w39[15]; //: TAP g64 @(1510,-11) /sn:0 /R:1 /w:[ 0 31 32 ] /ss:1
  assign w4 = w39[1]; //: TAP g6 @(239,-11) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  _GGNXOR2 #(6) g50 (.I0(w30), .I1(w35), .Z(w33));   //: @(1080,156) /sn:0 /R:3 /w:[ 1 1 1 ]
  assign w3 = w38[1]; //: TAP g7 @(243,53) /sn:0 /R:1 /w:[ 0 3 4 ] /ss:1
  assign w26 = w39[8]; //: TAP g35 @(904,-10) /sn:0 /R:1 /w:[ 0 17 18 ] /ss:1
  _GGNXOR2 #(6) g56 (.I0(w57), .I1(w50), .Z(w37));   //: @(1258,154) /sn:0 /R:3 /w:[ 1 1 1 ]
  assign w53 = w39[13]; //: TAP g58 @(1330,-12) /sn:0 /R:1 /w:[ 0 27 28 ] /ss:1
  //: LED g68 (w38) @(1651,21) /sn:0 /w:[ 33 ] /type:1
  //: IN g9 (EN) @(-12,-81) /sn:0 /w:[ 0 ]
  assign w18 = w38[6]; //: TAP g22 @(714,56) /sn:0 /R:1 /w:[ 0 13 14 ] /ss:1
  assign w22 = w39[7]; //: TAP g31 @(783,-10) /sn:0 /R:1 /w:[ 0 15 16 ] /ss:1
  //: LED g67 (w39) @(1609,-35) /sn:0 /w:[ 33 ] /type:1
  _GGNXOR2 #(6) g33 (.I0(w18), .I1(w23), .Z(w21));   //: @(708,152) /sn:0 /R:3 /w:[ 1 1 1 ]
  _GGNXOR2 #(6) g36 (.I0(w27), .I1(w28), .Z(w24));   //: @(972,157) /sn:0 /R:3 /w:[ 1 1 1 ]
  assign w28 = w39[9]; //: TAP g41 @(971,-10) /sn:0 /R:1 /w:[ 0 19 20 ] /ss:1
  _GGNXOR2 #(6) g45 (.I0(w29), .I1(w34), .Z(w32));   //: @(1152,158) /sn:0 /R:3 /w:[ 1 1 0 ]
  assign w54 = w38[15]; //: TAP g54 @(1514,59) /sn:0 /R:1 /w:[ 0 31 32 ] /ss:1
  //: OUT g42 (Out) @(682,418) /sn:0 /w:[ 1 ]
  assign w50 = w39[12]; //: TAP g52 @(1256,-12) /sn:0 /R:1 /w:[ 0 25 26 ] /ss:1
  _GGNXOR2 #(6) g66 (.I0(w56), .I1(w62), .Z(w59));   //: @(1438,155) /sn:0 /R:3 /w:[ 1 1 0 ]
  _GGNXOR2 #(6) g12 (.I0(w9), .I1(w10), .Z(w6));   //: @(421,155) /sn:0 /R:3 /w:[ 1 1 1 ]
  _GGNXOR2 #(6) g28 (.I0(w17), .I1(w22), .Z(w20));   //: @(780,154) /sn:0 /R:3 /w:[ 1 1 0 ]
  assign w31 = w38[8]; //: TAP g46 @(906,59) /sn:0 /R:1 /w:[ 0 17 18 ] /ss:1
  assign w0 = w38[0]; //: TAP g5 @(173,53) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  assign w8 = w39[2]; //: TAP g11 @(345,-10) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  assign w10 = w39[3]; //: TAP g14 @(422,-10) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  assign w14 = w39[4]; //: TAP g19 @(526,-10) /sn:0 /R:1 /w:[ 0 9 10 ] /ss:1
  assign w17 = w38[7]; //: TAP g21 @(784,56) /sn:0 /R:1 /w:[ 0 15 16 ] /ss:1
  _GGNXOR2 #(6) g61 (.I0(w54), .I1(w61), .Z(w58));   //: @(1510,157) /sn:0 /R:3 /w:[ 1 1 1 ]
  _GGNXOR2 #(6) g20 (.I0(w15), .I1(w16), .Z(w12));   //: @(600,153) /sn:0 /R:3 /w:[ 1 1 1 ]
  assign w62 = w39[14]; //: TAP g63 @(1436,-11) /sn:0 /R:1 /w:[ 0 29 30 ] /ss:1
  //: IN g0 (Reg1) @(60,-9) /sn:0 /w:[ 0 ]
  assign w30 = w38[10]; //: TAP g38 @(1086,60) /sn:0 /R:1 /w:[ 0 21 22 ] /ss:1
  _GGBUFIF16 #(4, 6) g15 (.Z(w38), .I(Reg2), .E(EN));   //: @(83,57) /sn:0 /w:[ 0 0 5 ]
  assign w15 = w38[5]; //: TAP g27 @(604,55) /sn:0 /R:1 /w:[ 0 11 12 ] /ss:1
  assign w34 = w39[11]; //: TAP g48 @(1152,-10) /sn:0 /R:1 /w:[ 0 23 24 ] /ss:1
  assign w29 = w38[11]; //: TAP g37 @(1156,60) /sn:0 /R:1 /w:[ 0 23 24 ] /ss:1
  assign w57 = w38[12]; //: TAP g62 @(1264,58) /sn:0 /R:1 /w:[ 0 25 26 ] /ss:1
  assign w56 = w38[14]; //: TAP g55 @(1444,59) /sn:0 /R:1 /w:[ 0 29 30 ] /ss:1
  _GGNXOR2 #(6) g13 (.I0(w11), .I1(w8), .Z(w7));   //: @(347,150) /sn:0 /R:3 /w:[ 1 1 0 ]
  _GGNXOR2 #(6) g53 (.I0(w52), .I1(w53), .Z(w36));   //: @(1330,156) /sn:0 /R:3 /w:[ 1 1 1 ]

endmodule
//: /netlistEnd

//: /netlistBegin Register_File
module Register_File(Addr1, Addr2, Write_Data, RW1, Data_out2, Data_out1, CLR, CLK);
//: interface  /sz:(291, 95) /bd:[ Ti0>Addr1[1:0](40/291) Ti1>Write_Data[15:0](149/291) Ti2>Addr2[1:0](251/291) Li0>CLK(26/95) Li1>RW1(69/95) Ri0>CLR(49/95) Bo0<Data_out1[15:0](70/291) Bo1<Data_out2[15:0](242/291) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input [1:0] Addr2;    //: /sn:0 {0}(680,547)(680,618)(100,618)(100,432)(#:47,432){1}
output [15:0] Data_out2;    //: /sn:0 {0}(#:693,524)(717,524)(717,524)(739,524){1}
input [15:0] Write_Data;    //: /sn:0 {0}(301,206)(301,192)(#:402,192){1}
//: {2}(404,190)(404,100){3}
//: {4}(404,96)(404,92)(231,92){5}
//: {6}(229,90)(229,39){7}
//: {8}(227,92)(224,92)(224,78)(210,78)(210,69)(#:47,69){9}
//: {10}(402,98)(301,98)(301,114){11}
//: {12}(404,194)(404,273){13}
//: {14}(#:402,275)(301,275)(301,300){15}
//: {16}(404,277)(404,359)(301,359)(#:301,397){17}
input CLR;    //: /sn:0 {0}(357,552)(357,523)(357,523)(357,493){1}
output [15:0] Data_out1;    //: /sn:0 {0}(#:692,315)(729,315){1}
input [1:0] Addr1;    //: /sn:0 {0}(#:47,199)(79,199)(79,199)(115,199){1}
//: {2}(119,199)(#:141,199){3}
//: {4}(117,201)(117,268)(116,268)(116,336){5}
input CLK;    //: /sn:0 {0}(249,552)(249,420)(250,420)(250,409){1}
//: {2}(252,407)(264,407){3}
//: {4}(250,405)(250,312){5}
//: {6}(252,310)(257,310)(257,310)(264,310){7}
//: {8}(250,308)(250,218){9}
//: {10}(252,216)(257,216)(257,216)(264,216){11}
//: {12}(250,214)(250,124)(264,124){13}
input RW1;    //: /sn:0 {0}(47,275)(98,275)(98,275)(152,275){1}
//: {2}(154,273)(154,221){3}
//: {4}(154,277)(154,344)(121,344){5}
wire w13;    //: /sn:0 {0}(340,402)(355,402){1}
//: {2}(357,400)(357,307){3}
//: {4}(357,303)(357,213){5}
//: {6}(357,209)(357,119)(340,119){7}
//: {8}(355,211)(340,211){9}
//: {10}(355,305)(340,305){11}
//: {12}(357,404)(357,477){13}
wire w25;    //: /sn:0 {0}(170,181)(236,181)(236,142)(352,142)(352,129)(340,129){1}
wire [15:0] w3;    //: /sn:0 {0}(#:301,418)(301,433)(498,433){1}
//: {2}(502,433)(590,433)(590,333)(601,333){3}
//: {4}(605,333)(663,333){5}
//: {6}(#:603,335)(603,542)(664,542){7}
//: {8}(500,431)(500,376){9}
wire [15:0] w0;    //: /sn:0 {0}(#:301,135)(301,167)(510,167){1}
//: {2}(514,167)(652,167)(652,295){3}
//: {4}(654,297)(663,297){5}
//: {6}(#:652,299)(652,506)(664,506){7}
//: {8}(512,165)(512,121){9}
wire w22;    //: /sn:0 {0}(170,217)(184,217)(184,382)(343,382)(343,412)(340,412){1}
wire w29;    //: /sn:0 {0}(170,193)(218,193)(218,243)(346,243)(346,221)(340,221){1}
wire [15:0] w12;    //: /sn:0 {0}(#:301,227)(301,249)(514,249){1}
//: {2}(518,249)(635,249)(635,307){3}
//: {4}(637,309)(663,309){5}
//: {6}(#:635,311)(635,518)(664,518){7}
//: {8}(516,247)(516,227)(515,227)(515,198){9}
wire [15:0] w10;    //: /sn:0 {0}(#:301,321)(301,334)(503,334){1}
//: {2}(507,334)(579,334)(579,321)(616,321){3}
//: {4}(620,321)(663,321){5}
//: {6}(#:618,323)(618,530)(664,530){7}
//: {8}(505,332)(#:505,322)(506,322)(506,288){9}
wire w23;    //: /sn:0 {0}(170,205)(198,205)(198,330)(352,330)(352,315)(340,315){1}
wire [1:0] w1;    //: /sn:0 {0}(#:116,352)(116,701)(800,701)(800,347)(679,347)(679,338){1}
//: enddecls

  //: IN g4 (Addr1) @(45,199) /sn:0 /w:[ 0 ]
  //: joint g8 (Addr1) @(117, 199) /w:[ 2 -1 1 4 ]
  //: IN g16 (Addr2) @(45,432) /sn:0 /w:[ 1 ]
  //: IN g3 (Write_Data) @(45,69) /sn:0 /w:[ 9 ]
  //: joint g26 (w0) @(652, 297) /w:[ 4 3 -1 6 ]
  //: joint g17 (w0) @(512, 167) /w:[ 2 8 1 -1 ]
  //: IN g2 (RW1) @(45,275) /sn:0 /w:[ 0 ]
  //: OUT g30 (Data_out2) @(736,524) /sn:0 /w:[ 1 ]
  //: joint g23 (w3) @(500, 433) /w:[ 2 8 1 -1 ]
  //: joint g39 (w13) @(357, 305) /w:[ -1 4 10 3 ]
  //: OUT g1 (Data_out1) @(726,315) /sn:0 /w:[ 1 ]
  //: LED g24 (Write_Data) @(229,32) /sn:0 /w:[ 7 ] /type:3
  //: joint g29 (w3) @(603, 333) /w:[ 4 -1 3 6 ]
  //: LED g18 (w12) @(515,191) /sn:0 /w:[ 9 ] /type:3
  _GGMUX4x16 #(12, 12) g25 (.I0(w3), .I1(w10), .I2(w12), .I3(w0), .S(Addr2), .Z(Data_out2));   //: @(680,524) /sn:0 /R:1 /w:[ 7 7 7 7 0 0 ] /ss:0 /do:0
  _GGNDECODER4 #(4, 4) g10 (.I(Addr1), .E(RW1), .Z0(w22), .Z1(w23), .Z2(w29), .Z3(w25));   //: @(154,199) /sn:0 /R:1 /w:[ 3 3 0 0 0 0 ] /ss:0 /do:0
  _GGREG16 #(10, 10, 20) r1 (.Q(w10), .D(Write_Data), .EN(w23), .CLR(w13), .CK(CLK));   //: @(301,310) /w:[ 0 15 1 11 7 ]
  //: joint g6 (Write_Data) @(404, 192) /w:[ -1 2 1 12 ]
  _GGBUFIF2 #(4, 6) g7 (.Z(w1), .I(Addr1), .E(~RW1));   //: @(116,342) /sn:0 /R:3 /w:[ 0 5 5 ]
  //: joint g9 (RW1) @(154, 275) /w:[ -1 2 1 4 ]
  //: LED g22 (w3) @(500,369) /sn:0 /w:[ 9 ] /type:3
  //: joint g31 (Write_Data) @(229, 92) /w:[ 5 6 8 -1 ]
  _GGREG16 #(10, 10, 20) r3 (.Q(w0), .D(Write_Data), .EN(w25), .CLR(w13), .CK(CLK));   //: @(301,124) /w:[ 0 11 1 7 13 ]
  //: IN g36 (CLR) @(357,554) /sn:0 /R:1 /w:[ 0 ]
  _GGMUX4x16 #(12, 12) g42 (.I0(w3), .I1(w10), .I2(w12), .I3(w0), .S(w1), .Z(Data_out1));   //: @(679,315) /sn:0 /R:1 /w:[ 5 5 5 5 1 0 ] /ss:0 /do:0
  //: joint g40 (w13) @(357, 211) /w:[ -1 6 8 5 ]
  _GGREG16 #(10, 10, 20) r0 (.Q(w3), .D(Write_Data), .EN(w22), .CLR(w13), .CK(CLK));   //: @(301,407) /w:[ 0 17 1 0 3 ]
  //: joint g12 (CLK) @(250, 310) /w:[ 6 8 -1 5 ]
  //: joint g28 (w10) @(618, 321) /w:[ 4 -1 3 6 ]
  //: joint g5 (Write_Data) @(404, 275) /w:[ -1 13 14 16 ]
  //: IN g11 (CLK) @(249,554) /sn:0 /R:1 /w:[ 0 ]
  //: joint g14 (CLK) @(250, 407) /w:[ 2 4 -1 1 ]
  //: joint g19 (w12) @(516, 249) /w:[ 2 8 1 -1 ]
  //: joint g21 (w10) @(505, 334) /w:[ 2 8 1 -1 ]
  //: LED g20 (w10) @(506,281) /sn:0 /w:[ 9 ] /type:3
  //: joint g38 (w13) @(357, 402) /w:[ -1 2 1 12 ]
  //: joint g0 (Write_Data) @(404, 98) /w:[ -1 4 10 3 ]
  //: LED g15 (w0) @(512,114) /sn:0 /w:[ 9 ] /type:3
  //: joint g27 (w12) @(635, 309) /w:[ 4 3 -1 6 ]
  _GGNBUF #(2) g37 (.I(CLR), .Z(w13));   //: @(357,487) /sn:0 /R:1 /w:[ 1 13 ]
  //: joint g13 (CLK) @(250, 216) /w:[ 10 12 -1 9 ]
  _GGREG16 #(10, 10, 20) r2 (.Q(w12), .D(Write_Data), .EN(w29), .CLR(w13), .CK(CLK));   //: @(301,216) /w:[ 0 0 1 9 11 ]

endmodule
//: /netlistEnd

//: /netlistBegin ALU
module ALU(OUT, MODE, IN2, IN1, EN, OF);
//: interface  /sz:(148, 53) /bd:[ Ti0>IN1[15:0](19/148) Ti1>IN2[15:0](124/148) Li0>EN(37/53) Ri0>MODE[1:0](37/53) Bo0<OUT[15:0](35/148) Bo1<OF(115/148) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
output OF;    //: /sn:0 {0}(34,162)(108,162){1}
output [15:0] OUT;    //: /sn:0 {0}(454,510)(#:454,451){1}
input [15:0] IN1;    //: /sn:0 {0}(#:214,98)(214,31)(255,31){1}
//: {2}(257,29)(257,-32){3}
//: {4}(259,-34)(356,-34){5}
//: {6}(360,-34)(435,-34)(435,98){7}
//: {8}(358,-32)(358,98){9}
//: {10}(255,-34)(#:147,-34){11}
//: {12}(257,33)(#:257,98){13}
input EN;    //: /sn:0 {0}(41,130)(103,130)(103,122){1}
input [15:0] IN2;    //: /sn:0 {0}(#:147,-17)(287,-17){1}
//: {2}(291,-17)(311,-17){3}
//: {4}(315,-17)(388,-17){5}
//: {6}(392,-17)(468,-17)(468,98){7}
//: {8}(390,-15)(390,98){9}
//: {10}(313,-15)(313,64){11}
//: {12}(289,-15)(289,98){13}
supply0 w17;    //: /sn:0 {0}(114,177)(172,177)(172,165)(129,165){1}
input [1:0] MODE;    //: /sn:0 {0}(#:38,100)(59,100){1}
//: {2}(63,100)(90,100){3}
//: {4}(#:61,102)(61,438)(431,438){5}
supply0 w15;    //: /sn:0 {0}(347,216)(347,178)(332,178)(332,192){1}
wire [15:0] w6;    //: /sn:0 {0}(#:358,114)(358,148){1}
wire w16;    //: /sn:0 {0}(329,213)(329,223)(310,223)(310,160)(297,160){1}
wire w13;    //: /sn:0 {0}(129,160)(249,160){1}
wire [15:0] w7;    //: /sn:0 {0}(#:435,114)(435,142)(434,142)(434,147){1}
wire w4;    //: /sn:0 {0}(473,106)(482,106)(482,125)(453,125){1}
//: {2}(451,123)(451,106)(440,106){3}
//: {4}(451,127)(451,137)(135,137)(135,94)(119,94){5}
wire w3;    //: /sn:0 {0}(395,106)(400,106)(400,123)(367,123){1}
//: {2}(365,121)(365,106)(363,106){3}
//: {4}(365,125)(365,131)(126,131)(126,106)(119,106){5}
wire [15:0] w0;    //: /sn:0 {0}(#:214,114)(214,128)(255,128){1}
//: {2}(257,126)(#:257,114){3}
//: {4}(257,130)(257,146){5}
wire [15:0] w12;    //: /sn:0 {0}(536,186)(536,213)(440,213)(#:440,176){1}
wire [15:0] w10;    //: /sn:0 {0}(448,422)(448,345)(374,345)(#:374,177){1}
wire [15:0] w1;    //: /sn:0 {0}(#:310,85)(310,126)(291,126){1}
//: {2}(289,124)(#:289,114){3}
//: {4}(289,128)(289,146){5}
wire [15:0] w8;    //: /sn:0 {0}(#:468,114)(468,139)(466,139)(466,147){1}
wire [15:0] w14;    //: /sn:0 {0}(460,422)(#:460,176){1}
wire w11;    //: /sn:0 {0}(119,82)(125,82)(125,50)(241,50){1}
//: {2}(245,50)(306,50){3}
//: {4}(310,50)(327,50)(327,192){5}
//: {6}(308,52)(308,64){7}
//: {8}(243,52)(243,106)(219,106){9}
wire w2;    //: /sn:0 {0}(262,106)(273,106)(273,116){1}
//: {2}(275,118)(305,118)(305,106)(294,106){3}
//: {4}(271,118)(119,118){5}
wire [15:0] w5;    //: /sn:0 {0}(#:273,175)(273,360)(276,360){1}
//: {2}(276,360)(472,360)(#:472,422){3}
//: {4}(274,362)(#:274,382)(436,382)(436,422){5}
wire [15:0] w9;    //: /sn:0 {0}(#:390,114)(390,148){1}
//: enddecls

  //: OUT g4 (OUT) @(454,507) /sn:0 /R:3 /w:[ 0 ]
  _GGBUFIF16 #(4, 6) g8 (.Z(w1), .I(IN2), .E(w2));   //: @(289,104) /sn:0 /R:3 /w:[ 3 13 3 ]
  _GGMUX4x16 #(12, 12) g16 (.I0(w5), .I1(w10), .I2(w14), .I3(w5), .S(MODE), .Z(OUT));   //: @(454,438) /sn:0 /w:[ 5 0 0 3 5 1 ] /ss:0 /do:0
  //: IN g3 (MODE) @(36,100) /sn:0 /w:[ 0 ]
  //: joint g26 (w1) @(289, 126) /w:[ 1 2 -1 4 ]
  _GGDIV16 #(492, 492) g17 (.A(w7), .B(w8), .Q(w14), .R(w12));   //: @(450,163) /sn:0 /w:[ 1 1 1 1 ]
  //: IN g2 (IN2) @(145,-17) /sn:0 /w:[ 0 ]
  //: joint g23 (IN2) @(289, -17) /w:[ 2 -1 1 12 ]
  //: joint g30 (MODE) @(61, 100) /w:[ 2 -1 1 4 ]
  //: joint g24 (IN1) @(257, -34) /w:[ 4 -1 10 3 ]
  //: IN g1 (IN1) @(145,-34) /sn:0 /w:[ 11 ]
  //: LED g29 (w12) @(536,179) /sn:0 /w:[ 0 ] /type:3
  _GGBUFIF16 #(4, 6) g18 (.Z(w8), .I(IN2), .E(w4));   //: @(468,104) /sn:0 /R:3 /w:[ 0 7 0 ]
  _GGXOR2x16 #(8) g25 (.I0(IN2), .I1({16{w11}}), .Z(w1));   //: @(310,75) /sn:0 /R:3 /w:[ 11 7 0 ]
  _GGMUL16 #(252) g10 (.A(w6), .B(w9), .P(w10));   //: @(374,164) /sn:0 /w:[ 1 1 1 ]
  _GGADD16 #(132, 134, 126, 128) g6 (.A(w0), .B(w1), .S(w5), .CI(w16), .CO(w13));   //: @(273,162) /sn:0 /w:[ 5 5 0 1 1 ]
  _GGBUFIF16 #(4, 6) g7 (.Z(w0), .I(IN1), .E(w2));   //: @(257,104) /sn:0 /R:3 /w:[ 3 13 0 ]
  //: joint g9 (w2) @(273, 118) /w:[ 2 1 4 -1 ]
  //: joint g35 (w11) @(308, 50) /w:[ 4 -1 3 6 ]
  _GGBUFIF16 #(4, 6) g31 (.Z(w0), .I(IN1), .E(w11));   //: @(214,104) /sn:0 /R:3 /w:[ 0 0 9 ]
  //: joint g22 (IN1) @(358, -34) /w:[ 6 -1 5 8 ]
  //: joint g33 (w0) @(257, 128) /w:[ -1 2 1 4 ]
  //: GROUND g36 (w15) @(347,222) /sn:0 /w:[ 0 ]
  _GGBUFIF16 #(4, 6) g12 (.Z(w9), .I(IN2), .E(w3));   //: @(390,104) /sn:0 /R:3 /w:[ 0 9 0 ]
  //: joint g34 (w11) @(243, 50) /w:[ 2 -1 1 8 ]
  //: joint g28 (w5) @(274, 360) /w:[ 2 -1 1 4 ]
  _GGDECODER4 #(6, 6) g5 (.I(MODE), .E(EN), .Z0(w2), .Z1(w3), .Z2(w4), .Z3(w11));   //: @(103,100) /sn:0 /R:1 /w:[ 3 1 5 5 5 0 ] /ss:0 /do:0
  _GGBUFIF16 #(4, 6) g11 (.Z(w6), .I(IN1), .E(w3));   //: @(358,104) /sn:0 /R:3 /w:[ 0 9 3 ]
  _GGOR2 #(6) g14 (.I0(w15), .I1(w11), .Z(w16));   //: @(329,203) /sn:0 /R:3 /w:[ 1 5 0 ]
  //: joint g21 (IN2) @(390, -17) /w:[ 6 -1 5 8 ]
  _GGBUFIF16 #(4, 6) g19 (.Z(w7), .I(IN1), .E(w4));   //: @(435,104) /sn:0 /R:3 /w:[ 0 7 3 ]
  //: joint g32 (IN1) @(257, 31) /w:[ -1 2 1 12 ]
  //: joint g20 (w4) @(451, 125) /w:[ 1 2 -1 4 ]
  //: IN g0 (EN) @(39,130) /sn:0 /w:[ 0 ]
  //: OUT g15 (OF) @(37,162) /sn:0 /R:2 /w:[ 0 ]
  _GGOR2 #(6) g38 (.I0(w17), .I1(w13), .Z(OF));   //: @(118,162) /sn:0 /R:2 /w:[ 1 0 1 ]
  //: joint g27 (IN2) @(313, -17) /w:[ 4 -1 3 10 ]
  //: GROUND g37 (w17) @(108,177) /sn:0 /R:3 /w:[ 0 ]
  //: joint g13 (w3) @(365, 123) /w:[ 1 2 -1 4 ]

endmodule
//: /netlistEnd

//: /netlistBegin jump_module
module jump_module(JNE_enable, offset_enable, Status_flag);
//: interface  /sz:(381, 80) /bd:[ Li0>JNE_enable(16/80) Li1>Status_flag(32/80) Ro0<offset_enable(16/80) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input JNE_enable;    //: {0}(478,183)(563,183)(46:563,199)(569,199){1}
output offset_enable;    //: {0}(590,202)(717,202)(717,225)(20:941,225){1}
input Status_flag;    //: /sn:0 {0}(502,276)(443,276)(443,245)(359,245)(359,243)(349,243){1}
wire w0;    //: /sn:0 {0}(518,276)(554,276)(554,204)(569,204){1}
//: enddecls

  //: IN g4 (JNE_enable) @(476,183) /sn:0 /w:[ 0 ]
  _GGNBUF #(2) g6 (.I(Status_flag), .Z(w0));   //: @(508,276) /sn:0 /w:[ 0 0 ]
  //: OUT g9 (offset_enable) @(938,225) /sn:0 /w:[ 1 ]
  //: IN g5 (Status_flag) @(347,243) /sn:0 /w:[ 1 ]
  _GGAND2 #(6) g0 (.I0(JNE_enable), .I1(w0), .Z(offset_enable));   //: @(580,202) /sn:0 /w:[ 1 1 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin Instruction_Fetch
module Instruction_Fetch(IR_OUT, EN, PC_in);
//: interface  /sz:(200, 56) /bd:[ Ti0>PC_in[7:0](90/200) Li0>EN(25/56) Bo0<IR_OUT[15:0](90/200) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input EN;    //: /sn:0 {0}(484,347)(484,311)(487,311)(487,273){1}
output [15:0] IR_OUT;    //: /sn:0 {0}(#:568,243)(537,243)(537,246)(#:504,246){1}
input [7:0] PC_in;    //: /sn:0 {0}(#:399,245)(435,245)(435,248)(469,248){1}
//: enddecls

  //: OUT g3 (IR_OUT) @(565,243) /sn:0 /w:[ 0 ]
  //: IN g2 (EN) @(484,349) /sn:0 /R:1 /w:[ 0 ]
  //: IN g1 (PC_in) @(397,245) /sn:0 /w:[ 0 ]
  _GGROM8x16 #(10, 30) g0 (.A(PC_in), .D(IR_OUT), .OE(~EN));   //: @(487,247) /sn:0 /w:[ 1 1 1 ] /mem:"/home/props/sumtillN.mem"

endmodule
//: /netlistEnd

//: /netlistBegin Instruction_Decode
module Instruction_Decode(RW1, IN2_User, ALU_EN, ALU_MODE, MemAddr2, EN, Reg1, Reg2, RR, HLT, Jmp_EN, Cmp_EN, Imm2, IR_IN);
//: interface  /sz:(463, 178) /bd:[ Li0>EN(135/178) Li1>IR_IN[15:0](34/178) To0<IN2_User(161/463) Bo0<MemAddr2[7:0](403/463) Bo1<Imm2[7:0](348/463) Bo2<Reg2[1:0](219/463) Bo3<Reg1[1:0](167/463) Bo4<ALU_EN(75/463) Bo5<ALU_MODE[1:0](29/463) Ro0<HLT(155/178) Ro1<RR(109/178) Ro2<Jmp_EN(77/178) Ro3<Cmp_EN(57/178) Ro4<RW1(27/178) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
output [7:0] Imm2;    //: /sn:0 {0}(#:708,243)(743,243){1}
output HLT;    //: /sn:0 {0}(421,279)(421,379)(573,379){1}
output [1:0] ALU_MODE;    //: /sn:0 {0}(#:266,369)(266,346)(230,346)(#:230,340){1}
output [1:0] Reg1;    //: /sn:0 {0}(#:526,330)(490,330)(#:490,167){1}
output IN2_User;    //: /sn:0 {0}(587,274)(587,309)(743,309){1}
input EN;    //: /sn:0 {0}(207,248)(304,248)(304,263)(326,263){1}
//: {2}(330,263)(371,263){3}
//: {4}(328,261)(328,241){5}
//: {6}(330,239)(535,239)(535,258)(545,258){7}
//: {8}(328,237)(328,141)(307,141)(307,158){9}
output Cmp_EN;    //: /sn:0 {0}(230,409)(230,396)(245,396)(245,441)(446,441)(446,431){1}
//: {2}(448,429)(512,429){3}
//: {4}(444,429)(415,429){5}
//: {6}(413,427)(413,340)(322,340)(322,354)(306,354){7}
//: {8}(411,429)(389,429)(389,279){9}
output [1:0] Reg2;    //: /sn:0 {0}(#:708,217)(740,217)(740,218)(743,218){1}
output Jmp_EN;    //: /sn:0 {0}(506,407)(393,407)(393,279){1}
input [15:0] IR_IN;    //: /sn:0 {0}(#:235,163)(299,163){1}
output [7:0] MemAddr2;    //: /sn:0 {0}(#:708,272)(743,272){1}
output ALU_EN;    //: /sn:0 {0}(511,500)(356,500)(356,364){1}
output RW1;    //: /sn:0 {0}(243,451)(659,451){1}
output RR;    //: /sn:0 {0}(330,434)(348,434)(348,572)(822,572)(822,187){1}
//: {2}(824,185)(863,185){3}
//: {4}(820,185)(694,185)(694,200){5}
//: {6}(696,202)(700,202)(700,212){7}
//: {8}(692,202)(637,202)(637,283)(551,283)(551,274){9}
wire [1:0] w6;    //: /sn:0 {0}(#:569,167)(569,245){1}
wire w16;    //: /sn:0 {0}(417,279)(417,294){1}
wire w13;    //: /sn:0 {0}(407,279)(407,294){1}
wire w7;    //: /sn:0 {0}(330,429)(346,429)(346,404)(366,404){1}
//: {2}(370,404)(386,404)(386,279){3}
//: {4}(368,406)(368,412)(371,412)(371,427){5}
wire w4;    //: /sn:0 {0}(361,343)(361,325)(315,325)(315,297)(375,297)(375,279){1}
wire [1:0] w22;    //: /sn:0 {0}(#:672,167)(672,217)(692,217){1}
wire [3:0] w0;    //: /sn:0 {0}(#:395,167)(395,232){1}
//: {2}(395,233)(395,250){3}
wire w3;    //: /sn:0 {0}(356,343)(356,328)(312,328)(312,293)(372,293)(372,279){1}
wire w20;    //: /sn:0 {0}(700,267)(700,254)(647,254)(647,301)(575,301)(575,274){1}
wire w18;    //: /sn:0 {0}(275,430)(275,422)(259,422)(259,406){1}
//: {2}(261,404)(300,404)(300,431)(309,431){3}
//: {4}(257,404)(240,404)(240,409){5}
wire w19;    //: /sn:0 {0}(700,238)(700,232)(642,232)(642,292)(563,292)(563,274){1}
wire w12;    //: /sn:0 {0}(403,279)(403,294){1}
wire w10;    //: /sn:0 {0}(396,279)(396,294){1}
wire w23;    //: /sn:0 {0}(235,430)(235,446){1}
wire w24;    //: /sn:0 {0}(290,354)(277,354)(277,340)(268,340)(268,332)(235,332){1}
wire [7:0] w21;    //: /sn:0 {0}(#:626,167)(626,241){1}
//: {2}(628,243)(692,243){3}
//: {4}(#:626,245)(626,272)(692,272){5}
wire [15:0] w1;    //: /sn:0 {0}(#:315,163)(394,163){1}
//: {2}(395,163)(489,163){3}
//: {4}(490,163)(568,163){5}
//: {6}(569,163)(625,163){7}
//: {8}(626,163)(671,163){9}
//: {10}(672,163)(775,163)(775,147){11}
wire w8;    //: /sn:0 {0}(189,435)(189,440)(220,440){1}
//: {2}(222,438)(222,390)(229,390){3}
//: {4}(233,390)(303,390)(303,389)(335,389){5}
//: {6}(339,389)(382,389)(382,279){7}
//: {8}(337,387)(337,379)(331,379)(331,331)(346,331)(346,343){9}
//: {10}(231,392)(231,401)(235,401)(235,409){11}
//: {12}(222,442)(222,451)(227,451){13}
wire w14;    //: /sn:0 {0}(410,279)(410,294){1}
wire w11;    //: /sn:0 {0}(400,279)(400,294){1}
wire w2;    //: /sn:0 {0}(351,343)(351,335)(308,335)(308,289)(368,289)(368,279){1}
wire w15;    //: /sn:0 {0}(414,279)(414,294){1}
wire w5;    //: /sn:0 {0}(366,343)(366,322)(319,322)(319,300)(379,300)(379,279){1}
wire [1:0] w9;    //: /sn:0 {0}(230,324)(230,312)(#:266,312)(266,298)(#:256,298)(256,233)(#:390,233){1}
//: enddecls

  //: OUT g8 (RW1) @(656,451) /sn:0 /w:[ 1 ]
  //: OUT g4 (IN2_User) @(740,309) /sn:0 /w:[ 1 ]
  //: joint g44 (w8) @(222, 440) /w:[ -1 2 1 12 ]
  //: joint g16 (EN) @(328, 263) /w:[ 2 4 1 -1 ]
  //: OUT g3 (ALU_EN) @(508,500) /sn:0 /w:[ 0 ]
  _GGBUFIF2 #(4, 6) g26 (.Z(Reg2), .I(w22), .E(RR));   //: @(698,217) /sn:0 /w:[ 0 1 7 ]
  _GGDECODER4 #(6, 6) g17 (.I(w6), .E(EN), .Z0(RR), .Z1(w19), .Z2(w20), .Z3(IN2_User));   //: @(569,258) /sn:0 /w:[ 1 7 9 1 1 0 ] /ss:0 /do:0
  //: OUT g2 (ALU_MODE) @(266,366) /sn:0 /R:3 /w:[ 0 ]
  //: OUT g23 (MemAddr2) @(740,272) /sn:0 /w:[ 1 ]
  _GGOR3 #(8) g30 (.I0(w18), .I1(w8), .I2(Cmp_EN), .Z(w23));   //: @(235,420) /sn:0 /R:3 /w:[ 5 11 0 0 ]
  _GGBUFIF8 #(4, 6) g24 (.Z(MemAddr2), .I(w21), .E(w20));   //: @(698,272) /sn:0 /w:[ 0 5 0 ]
  //: IN g1 (EN) @(205,248) /sn:0 /w:[ 0 ]
  //: joint g39 (RR) @(694, 202) /w:[ 6 5 8 -1 ]
  //: LED g29 (w1) @(775,140) /sn:0 /w:[ 11 ] /type:3
  assign w6 = w1[9:8]; //: TAP g18 @(569,161) /sn:0 /R:1 /w:[ 0 5 6 ] /ss:1
  //: joint g25 (w21) @(626, 243) /w:[ 2 1 -1 4 ]
  assign w0 = w1[15:12]; //: TAP g10 @(395,161) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:1
  //: OUT g6 (Reg1) @(523,330) /sn:0 /w:[ 0 ]
  _GGNBUF #(2) g35 (.I(Cmp_EN), .Z(w24));   //: @(300,354) /sn:0 /R:2 /w:[ 7 0 ]
  assign w21 = w1[7:0]; //: TAP g7 @(626,161) /sn:0 /R:1 /w:[ 0 7 8 ] /ss:1
  _GGDECODER16 #(6, 6) g9 (.I(w0), .E(EN), .Z0(w2), .Z1(w3), .Z2(w4), .Z3(w5), .Z4(w8), .Z5(w7), .Z6(Cmp_EN), .Z7(Jmp_EN), .Z8(w10), .Z9(w11), .Z10(w12), .Z11(w13), .Z12(w14), .Z13(w15), .Z14(w16), .Z15(HLT));   //: @(395,263) /sn:0 /w:[ 3 3 1 1 1 1 7 3 9 1 0 0 0 0 0 0 0 0 ] /ss:0 /do:0
  //: OUT g22 (Reg2) @(740,218) /sn:0 /w:[ 1 ]
  //: joint g31 (w8) @(231, 390) /w:[ 4 -1 3 10 ]
  //: joint g36 (Cmp_EN) @(446, 429) /w:[ 2 -1 4 1 ]
  //: LED g41 (w18) @(275,437) /sn:0 /R:2 /w:[ 0 ] /type:0
  //: LED g45 (w7) @(371,434) /sn:0 /R:2 /w:[ 5 ] /type:0
  _GGBUFIF2 #(4, 6) g33 (.Z(ALU_MODE), .I(w9), .E(w24));   //: @(230,330) /sn:0 /R:3 /w:[ 1 0 1 ]
  _GGOR2 #(6) g52 (.I0(RR), .I1(w7), .Z(w18));   //: @(319,431) /sn:0 /R:2 /w:[ 0 0 3 ]
  //: joint g42 (w7) @(368, 404) /w:[ 2 -1 1 4 ]
  //: OUT g40 (RR) @(860,185) /sn:0 /w:[ 3 ]
  assign w9 = w0[1:0]; //: TAP g12 @(393,233) /sn:0 /R:2 /w:[ 1 2 1 ] /ss:0
  //: OUT g46 (HLT) @(570,379) /sn:0 /w:[ 1 ]
  //: OUT g28 (Jmp_EN) @(503,407) /sn:0 /w:[ 0 ]
  //: joint g34 (Cmp_EN) @(413, 429) /w:[ 5 6 8 -1 ]
  _GGBUFIF16 #(4, 6) g14 (.Z(w1), .I(IR_IN), .E(EN));   //: @(305,163) /sn:0 /w:[ 0 1 9 ]
  _GGOR5 #(12) g11 (.I0(w5), .I1(w4), .I2(w3), .I3(w2), .I4(w8), .Z(ALU_EN));   //: @(356,354) /sn:0 /R:3 /w:[ 0 0 0 0 9 1 ]
  //: OUT g5 (Cmp_EN) @(509,429) /sn:0 /w:[ 3 ]
  //: OUT g21 (Imm2) @(740,243) /sn:0 /w:[ 1 ]
  //: joint g19 (EN) @(328, 239) /w:[ 6 8 -1 5 ]
  _GGBUFIF8 #(4, 6) g20 (.Z(Imm2), .I(w21), .E(w19));   //: @(698,243) /sn:0 /w:[ 0 3 0 ]
  //: joint g32 (w18) @(259, 404) /w:[ 2 -1 4 1 ]
  assign Reg1 = w1[11:10]; //: TAP g15 @(490,161) /sn:0 /R:1 /w:[ 1 3 4 ] /ss:1
  //: IN g0 (IR_IN) @(233,163) /sn:0 /w:[ 0 ]
  //: joint g38 (w8) @(337, 389) /w:[ 6 8 5 -1 ]
  //: LED g43 (w8) @(189,428) /sn:0 /w:[ 0 ] /type:0
  assign w22 = w1[7:6]; //: TAP g27 @(672,161) /sn:0 /R:1 /w:[ 0 9 10 ] /ss:1
  //: joint g37 (RR) @(822, 185) /w:[ 2 -1 4 1 ]
  _GGBUFIF #(4, 6) g13 (.Z(RW1), .I(w8), .E(w23));   //: @(233,451) /sn:0 /w:[ 0 13 1 ]

endmodule
//: /netlistEnd

//: /netlistBegin Control_Unit
module Control_Unit(OP_Forwarding, EN1, CLR, EN_Decoder, OP2, OP1, EN3, EN4, CLK, EN2);
//: interface  /sz:(250, 119) /bd:[ Ti0>OP2[1:0](166/250) Ti1>OP1[1:0](64/250) Li0>CLR(71/119) Li1>EN_Decoder(55/119) Li2>CLK(26/119) Bo0<EN4(190/250) Bo1<EN3(143/250) Bo2<EN2(95/250) Bo3<EN1(45/250) Ro0<OP_Forwarding(38/119) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
output EN3;    //: /sn:0 {0}(459,806)(343,806)(343,752){1}
supply0 w1;    //: /sn:0 {0}(369,514)(369,509)(423,509)(423,488)(351,488){1}
output EN4;    //: /sn:0 {0}(355,752)(355,818)(459,818){1}
input [1:0] OP1;    //: /sn:0 {0}(#:611,426)(611,384)(#:565,384){1}
input [1:0] OP2;    //: /sn:0 {0}(#:567,345)(698,345)(#:698,426){1}
input CLR;    //: /sn:0 {0}(473,516)(483,516)(483,560)(363,560){1}
input EN_Decoder;    //: /sn:0 {0}(280,736)(313,736){1}
input CLK;    //: /sn:0 {0}(252,565)(287,565){1}
output OP_Forwarding;    //: /sn:0 {0}(669,655)(655,655)(655,523){1}
output EN2;    //: /sn:0 {0}(331,752)(331,794)(459,794){1}
output EN1;    //: /sn:0 {0}(319,752)(319,783)(459,783){1}
reg [7:0] w5;    //: /sn:0 {0}(#:393,390)(393,399)(343,399)(343,474){1}
supply0 w9;    //: /sn:0 {0}(413,603)(413,570)(363,570){1}
wire w4;    //: /sn:0 {0}(243,480)(243,488)(303,488){1}
wire [1:0] w3;    //: /sn:0 {0}(#:337,723)(337,685){1}
wire [7:0] w0;    //: /sn:0 {0}(324,555)(#:324,503){1}
wire [7:0] w10;    //: /sn:0 {0}(#:311,474)(311,398)(189,398)(189,600)(322,600){1}
//: {2}(326,600)(347,600)(347,681)(337,681){3}
//: {4}(336,681)(180,681)(180,661){5}
//: {6}(324,598)(#:324,576){7}
//: enddecls

  //: OUT g8 (OP_Forwarding) @(666,655) /sn:0 /w:[ 0 ]
  //: OUT g4 (EN1) @(456,783) /sn:0 /w:[ 1 ]
  //: joint g3 (w10) @(324, 600) /w:[ 2 6 1 -1 ]
  //: IN g16 (CLR) @(471,516) /sn:0 /w:[ 0 ]
  //: IN g17 (EN_Decoder) @(278,736) /sn:0 /w:[ 0 ]
  //: IN g2 (OP2) @(565,345) /sn:0 /w:[ 0 ]
  //: LED g23 (w10) @(180,654) /sn:0 /w:[ 5 ] /type:1
  //: IN g1 (OP1) @(563,384) /sn:0 /w:[ 1 ]
  _GGREG8 #(10, 10, 20) g18 (.Q(w10), .D(w0), .EN(w9), .CLR(~CLR), .CK(CLK));   //: @(324,565) /sn:0 /w:[ 7 0 1 1 1 ]
  //: DIP g10 (w5) @(393,380) /sn:0 /w:[ 0 ] /st:1 /dn:1
  //: OUT g6 (EN3) @(456,806) /sn:0 /w:[ 0 ]
  _GGADD8 #(68, 70, 62, 64) g9 (.A(w10), .B(w5), .S(w0), .CI(w1), .CO(w4));   //: @(327,490) /sn:0 /w:[ 0 1 1 1 1 ]
  //: OUT g7 (EN4) @(456,818) /sn:0 /w:[ 1 ]
  //: IN g12 (CLK) @(250,565) /sn:0 /w:[ 0 ]
  //: GROUND g14 (w9) @(413,609) /sn:0 /w:[ 0 ]
  _GGDECODER4 #(6, 6) g11 (.I(w3), .E(EN_Decoder), .Z0(EN1), .Z1(EN2), .Z2(EN3), .Z3(EN4));   //: @(337,736) /sn:0 /w:[ 0 1 0 0 1 0 ] /ss:0 /do:0
  //: OUT g5 (EN2) @(456,794) /sn:0 /w:[ 1 ]
  assign w3 = w10[1:0]; //: TAP g21 @(337,679) /sn:0 /R:1 /w:[ 1 4 3 ] /ss:1
  Comparator_2bit g0 (.Reg1(OP1), .Reg2(OP2), .Out(OP_Forwarding));   //: @(593, 427) /sz:(133, 95) /sn:0 /p:[ Ti0>0 Ti1>1 Bo0<1 ]
  //: LED g15 (w4) @(243,473) /sn:0 /w:[ 0 ] /type:0
  //: GROUND g13 (w1) @(369,520) /sn:0 /w:[ 0 ]

endmodule
//: /netlistEnd

